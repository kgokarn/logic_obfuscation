module error_tolerant_type2_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339;

  xor U171 ( result_o[9], n143, add2_i[9]);
  xor U172 ( result_o[8], n144, add2_i[8]);
  xor U173 ( result_o[7], n145, n146);
  xor U174 ( n146, add2_i[7], add1_i[7]);
  xor U175 ( result_o[6], add2_i[6], n149);
  xor U176 ( n149, n150, add1_i[6]);
  xor U177 ( result_o[5], n153, add2_i[5]);
  xor U178 ( n153, n154, add1_i[5]);
  xor U179 ( result_o[4], n157, add2_i[4]);
  xor U180 ( n157, n158, add1_i[4]);
  xor U181 ( result_o[3], n171, n172);
  xor U182 ( n172, add2_i[3], add1_i[3]);
  xor U183 ( result_o[31], n188, n189);
  xor U184 ( n189, add2_i[31], add1_i[31]);
  xor U185 ( result_o[30], add2_i[30], n192);
  xor U186 ( n192, n193, add1_i[30]);
  xor U187 ( result_o[2], add2_i[2], n175);
  xor U188 ( n175, n176, add1_i[2]);
  xor U189 ( result_o[29], n196, add2_i[29]);
  xor U190 ( n196, n197, add1_i[29]);
  xor U191 ( result_o[28], n204, add2_i[28]);
  xor U192 ( n204, n205, add1_i[28]);
  xor U193 ( result_o[27], n217, n218);
  xor U194 ( n218, add2_i[27], add1_i[27]);
  xor U195 ( result_o[26], add2_i[26], n221);
  xor U196 ( n221, n222, add1_i[26]);
  xor U197 ( result_o[25], n225, add2_i[25]);
  xor U198 ( n225, n226, add1_i[25]);
  xor U199 ( result_o[24], n229, add2_i[24]);
  xor U200 ( n229, n230, add1_i[24]);
  xor U201 ( result_o[23], n242, n243);
  xor U202 ( n243, add2_i[23], add1_i[23]);
  xor U203 ( result_o[22], add2_i[22], n246);
  xor U204 ( n246, n247, add1_i[22]);
  xor U205 ( result_o[21], n250, add2_i[21]);
  xor U206 ( n250, n251, add1_i[21]);
  xor U207 ( result_o[20], n254, add2_i[20]);
  xor U208 ( n254, n255, add1_i[20]);
  xor U209 ( result_o[1], n201, add2_i[1]);
  xor U210 ( n201, n200, add1_i[1]);
  xor U211 ( result_o[19], n267, n268);
  xor U212 ( n268, add2_i[19], add1_i[19]);
  xor U213 ( result_o[18], add2_i[18], n271);
  xor U214 ( n271, n272, add1_i[18]);
  xor U215 ( result_o[17], n275, add2_i[17]);
  xor U216 ( n275, n276, add1_i[17]);
  xor U217 ( result_o[16], n279, add2_i[16]);
  xor U218 ( n279, n280, add1_i[16]);
  xor U219 ( result_o[15], n292, n293);
  xor U220 ( n293, add2_i[15], add1_i[15]);
  xor U221 ( result_o[14], add2_i[14], n296);
  xor U222 ( n296, n297, add1_i[14]);
  xor U223 ( result_o[13], n300, add2_i[13]);
  xor U224 ( n300, n301, add1_i[13]);
  xor U225 ( result_o[12], n304, add2_i[12]);
  xor U226 ( n304, n305, add1_i[12]);
  xor U227 ( result_o[11], n317, n318);
  xor U228 ( n318, add2_i[11], add1_i[11]);
  xor U229 ( result_o[10], n321, add2_i[10]);
  xor U230 ( n321, n322, add1_i[10]);
  xor U231 ( n143, n325, add1_i[9]);
  xor U232 ( n144, n328, add1_i[8]);
  not U233 ( n142, n170);
  nand U234 ( result_o[0], n170, n200);
  nand U235 ( n317, n319, n320);
  nand U236 ( n319, add1_i[10], n322);
  nand U237 ( n148, n149, add2_i[6]);
  nand U238 ( n295, n296, add2_i[14]);
  nand U239 ( n270, n271, add2_i[18]);
  nand U240 ( n245, n246, add2_i[22]);
  nand U241 ( n220, n221, add2_i[26]);
  nand U242 ( n191, n192, add2_i[30]);
  nand U243 ( n320, n321, add2_i[10]);
  nand U244 ( n170, add2_i[0], add1_i[0]);
  nand U245 ( n154, n155, n156);
  nand U246 ( n155, add1_i[4], n158);
  nand U247 ( n156, n157, add2_i[4]);
  nand U248 ( n301, n302, n303);
  nand U249 ( n302, add1_i[12], n305);
  nand U250 ( n303, n304, add2_i[12]);
  nand U251 ( n276, n277, n278);
  nand U252 ( n277, add1_i[16], n280);
  nand U253 ( n278, n279, add2_i[16]);
  nand U254 ( n251, n252, n253);
  nand U255 ( n252, add1_i[20], n255);
  nand U256 ( n253, n254, add2_i[20]);
  nand U257 ( n226, n227, n228);
  nand U258 ( n227, add1_i[24], n230);
  nand U259 ( n228, n229, add2_i[24]);
  nand U260 ( n197, n202, n203);
  nand U261 ( n202, add1_i[28], n205);
  nand U262 ( n203, n204, add2_i[28]);
  nand U263 ( n150, n151, n152);
  nand U264 ( n151, add1_i[5], n154);
  nand U265 ( n152, n153, add2_i[5]);
  nand U266 ( n297, n298, n299);
  nand U267 ( n298, add1_i[13], n301);
  nand U268 ( n299, n300, add2_i[13]);
  nand U269 ( n272, n273, n274);
  nand U270 ( n273, add1_i[17], n276);
  nand U271 ( n274, n275, add2_i[17]);
  nand U272 ( n247, n248, n249);
  nand U273 ( n248, add1_i[21], n251);
  nand U274 ( n249, n250, add2_i[21]);
  nand U275 ( n222, n223, n224);
  nand U276 ( n223, add1_i[25], n226);
  nand U277 ( n224, n225, add2_i[25]);
  nand U278 ( n193, n194, n195);
  nand U279 ( n194, add1_i[29], n197);
  nand U280 ( n195, n196, add2_i[29]);
  nand U281 ( n325, n326, n327);
  nand U282 ( n326, add1_i[8], n328);
  nand U283 ( n327, add2_i[8], n144);
  nand U284 ( n322, n323, n324);
  nand U285 ( n323, add1_i[9], n325);
  nand U286 ( n324, add2_i[9], n143);
  nand U287 ( n328, n329, n330);
  nand U288 ( n329, add1_i[7], n332);
  nand U289 ( n330, add2_i[7], n331);
  or U290 ( n331, n332, add1_i[7]);
  nand U291 ( n305, n306, n307);
  nand U292 ( n306, add1_i[11], n309);
  nand U293 ( n307, add2_i[11], n308);
  or U294 ( n308, n309, add1_i[11]);
  nand U295 ( n280, n281, n282);
  nand U296 ( n281, add1_i[15], n284);
  nand U297 ( n282, add2_i[15], n283);
  or U298 ( n283, n284, add1_i[15]);
  nand U299 ( n255, n256, n257);
  nand U300 ( n256, add1_i[19], n259);
  nand U301 ( n257, add2_i[19], n258);
  or U302 ( n258, n259, add1_i[19]);
  nand U303 ( n230, n231, n232);
  nand U304 ( n231, add1_i[23], n234);
  nand U305 ( n232, add2_i[23], n233);
  or U306 ( n233, n234, add1_i[23]);
  nand U307 ( n205, n206, n207);
  nand U308 ( n206, add1_i[27], n209);
  nand U309 ( n207, add2_i[27], n208);
  or U310 ( n208, n209, add1_i[27]);
  nand U311 ( n336, n337, n338);
  nand U312 ( n337, add2_i[5], add1_i[5]);
  nand U313 ( n338, add1_i[4], n339, add2_i[4]);
  or U314 ( n339, add2_i[5], add1_i[5]);
  nand U315 ( n313, n314, n315);
  nand U316 ( n314, add2_i[9], add1_i[9]);
  nand U317 ( n315, add1_i[8], n316, add2_i[8]);
  or U318 ( n316, add2_i[9], add1_i[9]);
  nand U319 ( n288, n289, n290);
  nand U320 ( n289, add2_i[13], add1_i[13]);
  nand U321 ( n290, add1_i[12], n291, add2_i[12]);
  or U322 ( n291, add2_i[13], add1_i[13]);
  nand U323 ( n263, n264, n265);
  nand U324 ( n264, add2_i[17], add1_i[17]);
  nand U325 ( n265, add1_i[16], n266, add2_i[16]);
  or U326 ( n266, add2_i[17], add1_i[17]);
  nand U327 ( n238, n239, n240);
  nand U328 ( n239, add2_i[21], add1_i[21]);
  nand U329 ( n240, add1_i[20], n241, add2_i[20]);
  or U330 ( n241, add2_i[21], add1_i[21]);
  nand U331 ( n213, n214, n215);
  nand U332 ( n214, add2_i[25], add1_i[25]);
  nand U333 ( n215, add1_i[24], n216, add2_i[24]);
  or U334 ( n216, add2_i[25], add1_i[25]);
  nand U335 ( n162, n163, n164);
  nand U336 ( n163, add1_i[2], n166);
  nand U337 ( n164, add2_i[2], n165);
  or U338 ( n165, n166, add1_i[2]);
  nand U339 ( n332, n333, n334);
  nand U340 ( n333, add1_i[6], n336);
  nand U341 ( n334, add2_i[6], n335);
  or U342 ( n335, n336, add1_i[6]);
  nand U343 ( n309, n310, n311);
  nand U344 ( n310, add1_i[10], n313);
  nand U345 ( n311, add2_i[10], n312);
  or U346 ( n312, n313, add1_i[10]);
  nand U347 ( n284, n285, n286);
  nand U348 ( n285, add1_i[14], n288);
  nand U349 ( n286, add2_i[14], n287);
  or U350 ( n287, n288, add1_i[14]);
  nand U351 ( n259, n260, n261);
  nand U352 ( n260, add1_i[18], n263);
  nand U353 ( n261, add2_i[18], n262);
  or U354 ( n262, n263, add1_i[18]);
  nand U355 ( n234, n235, n236);
  nand U356 ( n235, add1_i[22], n238);
  nand U357 ( n236, add2_i[22], n237);
  or U358 ( n237, n238, add1_i[22]);
  nand U359 ( n209, n210, n211);
  nand U360 ( n210, add1_i[26], n213);
  nand U361 ( n211, add2_i[26], n212);
  or U362 ( n212, n213, add1_i[26]);
  nand U363 ( n158, n159, n160);
  nand U364 ( n159, add1_i[3], n162);
  nand U365 ( n160, add2_i[3], n161);
  or U366 ( n161, n162, add1_i[3]);
  nand U367 ( n145, n147, n148);
  nand U368 ( n147, add1_i[6], n150);
  nand U369 ( n292, n294, n295);
  nand U370 ( n294, add1_i[14], n297);
  nand U371 ( n267, n269, n270);
  nand U372 ( n269, add1_i[18], n272);
  nand U373 ( n242, n244, n245);
  nand U374 ( n244, add1_i[22], n247);
  nand U375 ( n217, n219, n220);
  nand U376 ( n219, add1_i[26], n222);
  nand U377 ( n188, n190, n191);
  nand U378 ( n190, add1_i[30], n193);
  nand U379 ( n166, n167, n168);
  nand U380 ( n167, add1_i[1], n142);
  nand U381 ( n168, add2_i[1], n169);
  or U382 ( n169, add1_i[1], n142);
  or U383 ( n200, add2_i[0], add1_i[0]);
  nand U384 ( n171, n173, n174);
  nand U385 ( n173, add1_i[2], n176);
  nand U386 ( n174, n175, add2_i[2]);
  nand U387 ( n176, n198, n199);
  nand U388 ( n199, add1_i[1], n200);
  nand U389 ( n198, n201, add2_i[1]);
  nand U390 ( n184, n185, n186);
  nand U391 ( n185, add2_i[29], add1_i[29]);
  nand U392 ( n186, add1_i[28], n187, add2_i[28]);
  or U393 ( n187, add2_i[29], add1_i[29]);
  nand U394 ( n180, n181, n182);
  nand U395 ( n181, add1_i[30], n184);
  nand U396 ( n182, add2_i[30], n183);
  or U397 ( n183, n184, add1_i[30]);
  nand U398 ( result_o[32], n177, n178);
  nand U399 ( n177, add1_i[31], n180);
  nand U400 ( n178, add2_i[31], n179);
  or U401 ( n179, n180, add1_i[31]);
endmodule
