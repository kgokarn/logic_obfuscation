library verilog;
use verilog.vl_types.all;
entity broke_array_multiplier8_tb is
end broke_array_multiplier8_tb;
