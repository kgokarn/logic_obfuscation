module lower_part_or_carry_lookahead_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75;

  xor U63 ( result_o[9], n16, n17);
  xor U64 ( n17, add2_i[9], add1_i[9]);
  xor U65 ( result_o[8], n18, n19);
  xor U66 ( n19, add2_i[8], add1_i[8]);
  xor U67 ( result_o[7], n20, n21);
  xor U68 ( n21, add2_i[7], add1_i[7]);
  xor U69 ( result_o[6], n22, n23);
  xor U70 ( n23, add2_i[6], add1_i[6]);
  xor U71 ( result_o[5], n24, n25);
  xor U72 ( n25, add2_i[5], add1_i[5]);
  xor U73 ( result_o[4], n26, n27);
  xor U74 ( n27, add2_i[4], add1_i[4]);
  xor U75 (  result_o[15], n31, n32);
  xor U76 ( n32, add2_i[15], add1_i[15]);
  xor U77 ( result_o[14], n36, n37);
  xor U78 ( n37, add2_i[14], add1_i[14]);
  xor U79 ( result_o[13], n41, n42);
  xor U80 ( n42, add2_i[13], add1_i[13]);
  xor U81 ( result_o[12], n46, n47);
  xor U82 ( n47, add2_i[12], add1_i[12]);
  xor U83 ( result_o[11], n51, n52);
  xor U84 ( n52, add2_i[11], add1_i[11]);
  xor U85 ( result_o[10], n56, n57);
  xor U86 ( n57, add2_i[10], add1_i[10]);
  nand U87 ( result_o[3], n15, n14);
  nand U88 ( n24, n73, n74);
  nand U89 ( n73, add2_i[4], add1_i[4]);
  nand U90 ( n74, add1_i[3], n75, add2_i[3]);
  or U91 ( n75, add2_i[4], add1_i[4]);
  nand U92 ( n22, n70, n71);
  nand U93 ( n70, add1_i[5], n24);
  nand U94 ( n71, add2_i[5], n72);
  or U95 ( n72, n24, add1_i[5]);
  nand U96 ( n20, n67, n68);
  nand U97 ( n67, add1_i[6], n22);
  nand U98 ( n68, add2_i[6], n69);
  or U99 ( n69, n22, add1_i[6]);
  nand U100 ( n18, n64, n65);
  nand U101 ( n64, add1_i[7], n20);
  nand U102 ( n65, add2_i[7], n66);
  or U103 ( n66, n20, add1_i[7]);
  nand U104 ( n16, n61, n62);
  nand U105 ( n61, add1_i[8], n18);
  nand U106 ( n62, add2_i[8], n63);
  or U107 ( n63, n18, add1_i[8]);
  nand U108 ( n56, n58, n59);
  nand U109 ( n58, add1_i[9], n16);
  nand U110 ( n59, add2_i[9], n60);
  or U111 ( n60, n16, add1_i[9]);
  nand U112 ( n51, n53, n54);
  nand U113 ( n53, add1_i[10], n56);
  nand U114 ( n54, add2_i[10], n55);
  or U115 ( n55, n56, add1_i[10]);
  nand U116 ( n46, n48, n49);
  nand U117 ( n48, add1_i[11], n51);
  nand U118 ( n49, add2_i[11], n50);
  or U119 ( n50, n51, add1_i[11]);
  nand U120 ( n41, n43, n44);
  nand U121 ( n43, add1_i[12], n46);
  nand U122 ( n44, add2_i[12], n45);
  or U123 ( n45, n46, add1_i[12]);
  nand U124 ( n36, n38, n39);
  nand U125 ( n38, add1_i[13], n41);
  nand U126 ( n39, add2_i[13], n40);
  or U127 ( n40, n41, add1_i[13]);
  nand U128 ( n31, n33, n34);
  nand U129 ( n33, add1_i[14], n36);
  nand U130 ( n34, add2_i[14], n35);
  or U131 ( n35, n36, add1_i[14]);
  nand U132 ( result_o[16], n28, n29);
  nand U133 ( n28, add1_i[15], n31);
  nand U134 ( n29, add2_i[15], n30);
  or U135 ( n30, n31, add1_i[15]);
  nor U136 ( n26, n14, n15);
  not U137 ( n14, add1_i[3]);
  not U138 ( n15, add2_i[3]);
  or U139 ( result_o[0], add1_i[0], add2_i[0]);
  or U140 ( result_o[1], add1_i[1], add2_i[1]);
  or U141 ( result_o[2], add1_i[2], add2_i[2]);
endmodule
