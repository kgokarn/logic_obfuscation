module traditional_multiplier8 ( op1_i, op2_i, product_o );
  input [7:0] op1_i;
  input [7:0] op2_i;
  output [15:0] product_o;
  wire   n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472;

  xor U308 ( product_o[9], n142, n143);
  xor U309 ( n143, n144, n145);
  xor U310 ( product_o[8], n146, n147);
  xor U311 ( n146, n148, n149);
  xor U312 ( product_o[7], n150, n151);
  xor U313 ( product_o[6], n152, n153);
  xor U315 ( product_o[4], n157, n156);
  xor U316 ( product_o[2], n160, n161);
  xor U317 ( product_o[1], n162, n163);
  xor U319 ( product_o[13], n185, n178);
  xor U320 ( n182, n184, n183);
  xor U321 ( n183, n171, n172);
  xor U322 ( n185, n177, n176);
  xor U323 ( n218, n193, n194);
  xor U324 ( n188, n189, n223);
  xor U325 ( product_o[11], n207, n225);
  xor U326 ( n225, n205, n206);
  xor U327 ( n207, n210, n211);
  xor U328 ( n210, n212, n213);
  xor U329 ( n212, n216, n217);
  xor U330 ( product_o[10], n257, n231);
  xor U331 ( n234, n236, n237);
  xor U332 ( n236, n240, n241);
  xor U333 ( n257, n229, n230);
  xor U334 ( n142, n285, n286);
  xor U335 ( n147, n290, n291);
  xor U336 ( n156, n310, n311);
  xor U337 ( n311, n314, n315);
  xor U338 ( n309, n318, n317);
  xor U339 ( n313, n325, n326);
  xor U340 ( n153, n301, n300);
  xor U341 ( n300, n327, n328);
  xor U342 ( n326, n331, n332);
  xor U343 ( n314, n333, n336);
  xor U344 ( n331, n345, n346);
  xor U345 ( n151, n295, n294);
  xor U346 ( n294, n296, n297);
  xor U347 ( n297, n347, n348);
  xor U348 ( n328, n351, n352);
  xor U349 ( n345, n362, n358);
  xor U350 ( n352, n372, n373);
  xor U351 ( n348, n378, n379);
  xor U352 ( n373, n388, n389);
  xor U353 ( n379, n396, n397);
  xor U354 ( n291, n398, n399);
  xor U355 ( n399, n408, n409);
  xor U356 ( n409, n414, n415);
  xor U357 ( n396, n422, n423);
  xor U358 ( n415, n432, n433);
  xor U359 ( n285, n434, n435);
  xor U360 ( n434, n260, n261);
  xor U361 ( n262, n270, n271);
  xor U362 ( n432, n449, n450);
  nand U364 ( n148, n151, n150);
  nand U365 ( n206, n226, n227);
  or U366 ( n226, n231, n230);
  nand U367 ( n227, n228, n229);
  nand U368 ( n228, n230, n231);
  and U369 ( n230, n282, n283);
  nand U370 ( n282, n145, n144);
  nand U371 ( n283, n142, n284);
  or U372 ( n284, n145, n144);
  nand U373 ( n144, n287, n288);
  or U374 ( n287, n148, n149);
  nand U375 ( n288, n147, n289);
  nand U376 ( n289, n149, n148);
  nand U377 ( n168, n173, n174);
  or U378 ( n173, n178, n177);
  nand U379 ( n174, n175, n176);
  nand U380 ( n175, n177, n178);
  and U381 ( n199, n202, n203);
  nand U382 ( n202, n207, n206);
  nand U383 ( n203, n204, n205);
  or U384 ( n204, n206, n207);
  xnor U385 ( n231, n234, n235);
  xnor U386 ( n155, n312, n313);
  nand U387 ( n312, n311, n310);
  xnor U388 ( n261, n263, n262);
  xnor U389 ( product_o[12], n200, n201);
  xnor U390 ( n201, n198, n199);
  nand U391 ( n152, n302, n303);
  nand U392 ( n302, n313, n310, n311);
  nand U393 ( n303, n155, n156, n157);
  nand U394 ( n145, n374, n375);
  nand U395 ( n374, n399, n398);
  nand U396 ( n375, n291, n290);
  and U397 ( n149, n292, n293);
  nand U398 ( n292, n296, n297);
  nand U399 ( n293, n294, n295);
  nand U400 ( n150, n298, n299);
  nand U401 ( n299, n300, n301);
  nand U402 ( n298, n153, n152);
  nand U403 ( n301, n329, n330);
  nand U404 ( n329, n331, n332);
  nand U405 ( n330, n325, n326);
  and U406 ( n177, n195, n196);
  or U407 ( n195, n200, n199);
  nand U408 ( n196, n197, n198);
  nand U409 ( n197, n199, n200);
  xnor U410 ( n178, n181, n182);
  nand U411 ( n198, n208, n209);
  nand U412 ( n208, n212, n213);
  nand U413 ( n209, n210, n211);
  xnor U414 ( product_o[5], n468, n155);
  nand U415 ( n468, n156, n157);
  nand U416 ( n176, n191, n192);
  nand U417 ( n192, n193, n194);
  nand U418 ( n205, n232, n233);
  nand U419 ( n232, n236, n237);
  nand U420 ( n233, n234, n235);
  nand U421 ( n229, n410, n411);
  nand U422 ( n410, n434, n435);
  nand U423 ( n411, n285, n286);
  nor U424 ( n296, n138, n354, n136);
  nor U425 ( n336, n140, n136);
  xnor U426 ( n395, n428, n429);
  nor U427 ( n429, n125, n141);
  xnor U428 ( n320, n341, n342);
  nor U429 ( n342, n133, n141);
  xnor U430 ( n344, n368, n369);
  nor U431 ( n369, n130, n141);
  xnor U432 ( n371, n392, n393);
  nor U433 ( n393, n127, n141);
  xnor U434 ( n305, n323, n324);
  nor U435 ( n324, n134, n141);
  xnor U436 ( n387, n406, n407);
  nor U437 ( n407, n140, n134);
  xnor U438 ( n431, n455, n456);
  nor U439 ( n456, n141, n124);
  xnor U440 ( n280, n281, n445);
  nor U441 ( n445, n140, n127);
  xnor U442 ( n358, n359, n363);
  nor U443 ( n363, n140, n135);
  xnor U444 ( n433, n451, n452);
  xnor U445 ( n315, n337, n338);
  xnor U446 ( n346, n364, n365);
  xnor U447 ( n397, n424, n425);
  xnor U448 ( n423, n442, n443);
  nor U449 ( n443, n133, n140);
  xnor U450 ( n450, n466, n467);
  nor U451 ( n467, n130, n140);
  nand U452 ( n310, n306, n316);
  nand U453 ( n316, n317, n318);
  nand U454 ( n263, n447, n448);
  nand U455 ( n447, n452, n451);
  or U456 ( n448, n433, n432);
  xnor U457 ( product_o[14], n469, n166);
  nor U458 ( n469, n167, n168);
  nand U459 ( n332, n334, n335);
  nand U460 ( n334, n338, n337);
  or U461 ( n335, n315, n314);
  nand U462 ( n378, n384, n385);
  nand U463 ( n384, n389, n388);
  nand U464 ( n385, n373, n372);
  nand U465 ( n295, n349, n350);
  nand U466 ( n349, n352, n351);
  nand U467 ( n350, n327, n328);
  nand U468 ( n290, n376, n377);
  nand U469 ( n376, n379, n378);
  nand U470 ( n377, n347, n348);
  nand U471 ( n398, n400, n380);
  nand U472 ( n351, n360, n361);
  nand U473 ( n360, n365, n364);
  or U474 ( n361, n346, n345);
  nand U475 ( n414, n420, n421);
  nand U476 ( n420, n425, n424);
  or U477 ( n421, n397, n396);
  and U478 ( n157, n158, n161, n160);
  or U479 ( n265, n137, n134, n460);
  or U480 ( n245, n137, n133, n274);
  or U481 ( n380, n136, n137, n383);
  or U482 ( n416, n137, n135, n419);
  nand U483 ( product_o[15], n164, n165);
  nand U484 ( n165, n166, n167);
  nand U485 ( n164, n166, n168);
  nor U486 ( n223, n138, n125);
  nor U487 ( n160, n141, n135, n162);
  nor U488 ( n181, n139, n190, n124);
  nor U489 ( n325, n333, n140, n136);
  nor U490 ( n189, n125, n139, n224);
  xnor U491 ( n217, n224, n246);
  nor U492 ( n246, n139, n125);
  xnor U493 ( n255, n256, n267);
  nor U494 ( n267, n140, n125);
  xnor U495 ( n190, n188, n222);
  nor U496 ( n222, n137, n127);
  xnor U497 ( n193, n190, n221);
  nor U498 ( n221, n139, n124);
  nor U499 ( n172, n124, n138);
  xnor U500 ( n241, n243, n242);
  nor U501 ( n171, n125, n137);
  nand U502 ( n191, n218, n217, n216);
  nand U503 ( n200, n191, n214);
  nand U504 ( n214, n122, n215);
  nand U505 ( n215, n216, n217);
  not U506 ( n122, n218);
  nand U507 ( n235, n258, n259);
  nand U508 ( n258, n262, n263);
  or U509 ( n259, n260, n261);
  nand U510 ( n237, n264, n265);
  nand U511 ( n213, n244, n245);
  nand U512 ( n435, n436, n416);
  nand U513 ( n194, n219, n220);
  nand U514 ( n211, n238, n239);
  nand U515 ( n238, n242, n243);
  or U516 ( n239, n240, n241);
  nand U517 ( n167, n179, n180);
  nand U518 ( n179, n183, n184);
  nand U519 ( n180, n181, n182);
  nand U520 ( n286, n412, n413);
  nand U521 ( n412, n415, n414);
  nand U522 ( n413, n408, n409);
  xnor U523 ( product_o[3], n158, n159);
  nand U524 ( n159, n160, n161);
  or U525 ( n220, n137, n130, n249);
  nand U526 ( n243, n268, n269);
  nand U527 ( n268, n270, n271);
  nor U528 ( product_o[0], n141, n136);
  xnor U529 ( n452, n446, n470);
  nand U530 ( n470, op1_i[6], op2_i[2]);
  not U531 ( n125, op1_i[6]);
  nand U532 ( n362, op1_i[0], op2_i[5]);
  nand U533 ( n422, op2_i[5], op1_i[2]);
  nand U534 ( n449, op2_i[5], op1_i[3]);
  xnor U535 ( n161, n304, n305);
  nand U536 ( n304, op1_i[0], op2_i[2]);
  not U537 ( n141, op2_i[0]);
  not U538 ( n140, op2_i[4]);
  xnor U539 ( n338, n343, n344);
  nand U540 ( n343, op2_i[2], op1_i[2]);
  xnor U541 ( n365, n370, n371);
  nand U542 ( n370, op2_i[2], op1_i[3]);
  xnor U543 ( n425, n430, n431);
  nand U544 ( n430, op2_i[2], op1_i[5]);
  xnor U545 ( n372, n386, n387);
  nand U546 ( n386, op1_i[1], op2_i[5]);
  not U547 ( n134, op1_i[2]);
  not U548 ( n133, op1_i[3]);
  not U549 ( n130, op1_i[4]);
  not U550 ( n127, op1_i[5]);
  not U551 ( n124, op1_i[7]);
  not U552 ( n136, op1_i[0]);
  xnor U553 ( n317, n319, n320);
  nand U554 ( n319, op2_i[2], op1_i[1]);
  xnor U555 ( n389, n394, n395);
  nand U556 ( n394, op2_i[2], op1_i[4]);
  nor U557 ( n327, n296, n353);
  and U558 ( n353, n354, n355);
  nand U559 ( n355, op1_i[0], op2_i[6]);
  not U560 ( n135, op1_i[1]);
  nand U561 ( n306, op1_i[0], op2_i[3], n309);
  nand U562 ( n400, op2_i[6], n403, op1_i[1]);
  nand U563 ( n436, op1_i[2], n439, op2_i[6]);
  nand U564 ( n264, op1_i[3], n463, op2_i[6]);
  nand U565 ( n337, n339, n340);
  or U566 ( n339, n141, n133, n341);
  nand U567 ( n340, op1_i[1], n320, op2_i[2]);
  nand U568 ( n341, op2_i[1], op1_i[2]);
  nand U569 ( n368, op2_i[1], op1_i[3]);
  nand U570 ( n392, op2_i[1], op1_i[4]);
  nand U571 ( n323, op2_i[1], op1_i[1]);
  nand U572 ( n406, op1_i[3], op2_i[3]);
  nand U573 ( n359, op1_i[2], op2_i[3]);
  nand U574 ( n428, op2_i[1], op1_i[5]);
  nand U575 ( n442, op2_i[3], op1_i[4]);
  nand U576 ( n455, op1_i[6], op2_i[1]);
  nand U577 ( n466, op1_i[5], op2_i[3]);
  nand U578 ( n383, n400, n401);
  nand U579 ( n401, n131, n402);
  nand U580 ( n402, op1_i[1], op2_i[6]);
  not U581 ( n131, n403);
  nand U582 ( n274, n244, n275);
  nand U583 ( n275, n126, n276);
  nand U584 ( n276, op2_i[6], op1_i[4]);
  not U585 ( n126, n277);
  and U586 ( n158, n306, n307);
  nand U587 ( n307, n132, n308);
  nand U588 ( n308, op1_i[0], op2_i[3]);
  not U589 ( n132, n309);
  nand U590 ( n424, n426, n427);
  or U591 ( n426, n141, n125, n428);
  nand U592 ( n427, op1_i[4], n395, op2_i[2]);
  nand U593 ( n364, n366, n367);
  or U594 ( n366, n141, n130, n368);
  nand U595 ( n367, op1_i[2], n344, op2_i[2]);
  nand U596 ( n318, n321, n322);
  or U597 ( n321, n141, n134, n323);
  nand U598 ( n322, op2_i[2], n305, op1_i[0]);
  nand U599 ( n388, n390, n391);
  or U600 ( n390, n141, n127, n392);
  nand U601 ( n391, op1_i[3], n371, op2_i[2]);
  nand U602 ( n403, n404, n405);
  or U603 ( n404, n134, n140, n406);
  nand U604 ( n405, op2_i[5], n387, op1_i[1]);
  nand U605 ( n451, n453, n454);
  or U606 ( n453, n124, n141, n455);
  nand U607 ( n454, op1_i[5], n431, op2_i[2]);
  nand U608 ( n277, n278, n279);
  or U609 ( n278, n127, n140, n281);
  nand U610 ( n279, op1_i[4], n280, op2_i[5]);
  nand U611 ( n333, op1_i[1], op2_i[3]);
  nand U612 ( n439, n440, n441);
  or U613 ( n440, n140, n133, n442);
  nand U614 ( n441, op1_i[2], n423, op2_i[5]);
  nand U615 ( n463, n464, n465);
  or U616 ( n464, n140, n130, n466);
  nand U617 ( n465, op1_i[3], n450, op2_i[5]);
  and U618 ( n446, op1_i[7], op2_i[1]);
  and U619 ( n347, n380, n381);
  nand U620 ( n381, n382, n383);
  nand U621 ( n382, op1_i[0], op2_i[7]);
  and U622 ( n408, n416, n417);
  nand U623 ( n417, n418, n419);
  nand U624 ( n418, op2_i[7], op1_i[1]);
  nand U625 ( n260, n265, n458);
  nand U626 ( n458, n459, n460);
  nand U627 ( n459, op2_i[7], op1_i[2]);
  nand U628 ( n240, n245, n272);
  nand U629 ( n272, n273, n274);
  nand U630 ( n273, op2_i[7], op1_i[3]);
  nor U631 ( n354, n471, n472);
  nor U632 ( n471, n135, n140, n359);
  and U633 ( n472, op2_i[5], n358, op1_i[0]);
  nand U634 ( n419, n436, n437);
  nand U635 ( n437, n129, n438);
  nand U636 ( n438, op2_i[6], op1_i[2]);
  not U637 ( n129, n439);
  nand U638 ( n460, n264, n461);
  nand U639 ( n461, n128, n462);
  nand U640 ( n462, op2_i[6], op1_i[3]);
  not U641 ( n128, n463);
  not U642 ( n137, op2_i[7]);
  xnor U643 ( n242, n266, n255);
  nand U644 ( n266, op1_i[5], op2_i[5]);
  xnor U645 ( n271, n444, n280);
  nand U646 ( n444, op2_i[5], op1_i[4]);
  not U647 ( n139, op2_i[5]);
  nand U648 ( n269, op2_i[2], op1_i[6], n446);
  not U649 ( n138, op2_i[6]);
  and U650 ( n216, n220, n247);
  nand U651 ( n247, n248, n249);
  nand U652 ( n248, op2_i[7], op1_i[4]);
  nand U653 ( n244, op1_i[4], n277, op2_i[6]);
  nand U654 ( n219, op2_i[6], n252, op1_i[5]);
  nand U655 ( n224, op1_i[7], op2_i[4]);
  nand U656 ( n281, op1_i[6], op2_i[3]);
  nand U657 ( n256, op1_i[7], op2_i[3]);
  nand U658 ( n249, n219, n250);
  nand U659 ( n250, n123, n251);
  nand U660 ( n251, op1_i[5], op2_i[6]);
  not U661 ( n123, n252);
  nand U662 ( n184, n186, n187);
  nand U663 ( n186, n189, op2_i[6]);
  nand U664 ( n187, op2_i[7], n188, op1_i[5]);
  nand U665 ( n252, n253, n254);
  or U666 ( n253, n125, n140, n256);
  nand U667 ( n254, op2_i[5], n255, op1_i[5]);
  nand U668 ( n162, op1_i[0], op2_i[1]);
  and U669 ( n270, op2_i[2], n269, op1_i[7]);
  nand U670 ( n163, op2_i[0], op1_i[1]);
  and U671 ( n166, op2_i[7], n170, op1_i[7]);
  nand U672 ( n170, n171, n172);
endmodule
