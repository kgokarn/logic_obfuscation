library verilog;
use verilog.vl_types.all;
entity error_tolerant_type2_adder16_tb is
end error_tolerant_type2_adder16_tb;
