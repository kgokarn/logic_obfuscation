library verilog;
use verilog.vl_types.all;
entity carry_lookahead_adder16_tb is
end carry_lookahead_adder16_tb;
