library verilog;
use verilog.vl_types.all;
entity traditional_multiplier8_tb is
end traditional_multiplier8_tb;
