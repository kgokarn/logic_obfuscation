module xnor_based_ripple_carry_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n178, n179, n180, n181, n183, n186, n187, n188, n189, n190, n191,
         n192, n193, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369;

  xor U138 ( result_o[8], add2_i[8], n345);
  xor U139 ( n203, add2_i[3], add1_i[3]);
  xor U144 ( result_o[29], add2_i[29], n331);
  xor U146 ( result_o[28], n227, n228);
  xor U149 ( result_o[25], n237, add2_i[25]);
  xor U151 ( result_o[24], n347, add2_i[24]);
  xor U153 ( result_o[22], add2_i[22], n250);
  xor U163 ( result_o[16], add2_i[16], n280);
  xor U165 ( result_o[15], n284, add2_i[15]);
  xor U167 ( result_o[14], add2_i[14], n288);
  xor U169 ( result_o[13], add2_i[13], n292);
  xor U171 ( result_o[12], add2_i[12], n296);
  xor U175 ( result_o[10], add2_i[10], n304);
  xor U177 ( n190, add1_i[7], add2_i[7]);
  xor U179 ( n199, add1_i[4], add2_i[4]);
  xor U180 ( n216, add1_i[2], add2_i[2]);
  xor U181 ( n267, add1_i[0], add2_i[0]);
  xnor U182 ( n326, n277, n348);
  not U183 ( n327, n210);
  not U184 ( n328, n327);
  or U185 ( n325, n217, n359, n218);
  nand U186 ( n340, n329, add1_i[18]);
  not U187 ( n329, n274);
  nand U188 ( n322, n183, n199, n201);
  nand U189 ( n339, n326, add2_i[17], add1_i[18]);
  nand U190 ( n313, n179, n321, n322, n315);
  and U191 ( n335, n339, add2_i[18], n340);
  nand U192 ( n320, n195, add2_i[5], add1_i[5]);
  nand U193 ( n249, n248, n251, add2_i[22]);
  xor U194 ( result_o[9], add2_i[9], n187);
  xor U195 ( result_o[11], add2_i[11], n300);
  xor U196 ( result_o[17], add2_i[17], n326);
  xor U197 ( result_o[19], add2_i[19], n263);
  xor U198 ( result_o[20], add2_i[20], n260);
  xor U199 ( result_o[21], add2_i[21], n255);
  xor U200 ( result_o[26], add2_i[26], n233);
  xor U201 ( result_o[30], add2_i[30], n328);
  xor U202 ( result_o[31], n206, add2_i[31]);
  not U203 ( n343, add1_i[24]);
  not U204 ( n342, add1_i[19]);
  not U205 ( n346, add1_i[25]);
  not U206 ( n330, n214);
  not U207 ( n331, n330);
  and U208 ( n332, n321, n322);
  nand U209 ( n333, n209, n208);
  and U210 ( n268, add1_i[1], add2_i[1]);
  or U211 ( n334, add1_i[0], add2_i[0]);
  nand U212 ( n270, n336, n335);
  or U213 ( n336, n273, add1_i[18]);
  nand U214 ( n337, n212, n213);
  nand U215 ( n338, n235, n236);
  and U216 ( n269, n339, n340);
  nand U217 ( n341, n231, n232);
  xnor U218 ( n263, n264, n342);
  xnor U219 ( n241, n242, n343);
  not U220 ( n344, n188);
  not U221 ( n345, n344);
  xnor U222 ( n237, n238, n346);
  not U223 ( n350, add1_i[13]);
  nor U224 ( n217, n334, n268);
  xor U225 ( n347, n242, add1_i[24]);
  not U226 ( n349, add1_i[15]);
  not U227 ( n348, add1_i[17]);
  xnor U228 ( n276, n277, n348);
  xnor U229 ( n284, n285, n349);
  xnor U230 ( n292, n293, n350);
  not U231 ( n351, add1_i[14]);
  not U232 ( n352, add1_i[16]);
  xnor U233 ( n288, n289, n351);
  xnor U234 ( n280, n281, n352);
  nor U235 ( n353, add1_i[0], add2_i[0], n367);
  not U236 ( n362, add1_i[29]);
  not U237 ( n355, add1_i[12]);
  not U238 ( n354, add1_i[20]);
  not U239 ( n356, add1_i[30]);
  xnor U240 ( n260, n259, n354);
  xnor U241 ( n296, n297, n355);
  xnor U242 ( n210, n211, n356);
  xor U243 ( n357, add1_i[6], add2_i[6]);
  not U244 ( n361, add1_i[21]);
  not U245 ( n358, add1_i[26]);
  not U246 ( n360, add1_i[31]);
  xnor U247 ( n233, n234, n358);
  xnor U248 ( n359, add1_i[2], add2_i[2]);
  xnor U249 ( n206, n207, n360);
  xnor U250 ( n255, n256, n361);
  xnor U251 ( n214, n215, n362);
  not U252 ( n183, n200);
  not U253 ( n181, n193);
  nor U254 ( result_o[7], n189, n190);
  nor U255 ( n189, n191, n192);
  nor U256 ( result_o[4], n199, n369, n200);
  not U257 ( result_o[0], n267);
  not U258 ( n366, add1_i[11]);
  not U259 ( n365, add1_i[9]);
  xor U260 ( n195, add1_i[6], add2_i[6]);
  xnor U261 ( n193, add1_i[5], add2_i[5]);
  nor U262 ( n218, add2_i[1], add1_i[1]);
  nor U263 ( n200, add2_i[3], add1_i[3]);
  nand U264 ( n319, add1_i[6], add2_i[6]);
  nand U265 ( n221, n222, n178);
  xnor U266 ( n228, add2_i[28], n178);
  xor U267 ( result_o[23], n363, n246);
  xor U268 ( n363, add1_i[23], add2_i[23]);
  and U269 ( n250, n251, n248);
  nand U270 ( n315, add2_i[7], add1_i[7]);
  nand U271 ( n321, add1_i[4], add2_i[4]);
  xnor U272 ( result_o[18], add2_i[18], n364);
  nand U273 ( n364, n269, n272);
  not U274 ( n178, add1_i[28]);
  not U275 ( n186, add2_i[27]);
  nor U276 ( n196, n197, n198);
  and U277 ( n198, add1_i[5], add2_i[5]);
  nor U278 ( result_o[1], n265, n266);
  nor U279 ( n265, n367, n218);
  nor U280 ( n266, add1_i[0], n267);
  and U281 ( n304, n305, n302);
  nand U282 ( n239, add1_i[24], n242);
  nand U283 ( n309, n310, n311);
  xnor U284 ( n187, n309, n365);
  xnor U285 ( n300, n366, n301);
  and U286 ( n367, add1_i[1], add2_i[1]);
  nand U287 ( n312, n315, n316);
  not U288 ( n179, n192);
  nand U289 ( n316, n190, n317);
  nand U290 ( n317, n179, n318);
  and U291 ( n368, n324, n323);
  and U292 ( n369, n202, n323);
  nand U293 ( n324, add1_i[2], add2_i[2]);
  nand U294 ( n323, add2_i[3], add1_i[3]);
  and U295 ( n202, n325, n324);
  nor U296 ( result_o[3], n202, n203);
  nand U297 ( n201, n325, n368);
  nand U298 ( n212, add1_i[29], n215);
  nand U299 ( n290, n293, add1_i[13]);
  nand U300 ( n298, add1_i[11], n301);
  nand U301 ( n307, n309, add1_i[9]);
  nand U302 ( n215, n219, n220);
  nand U303 ( n220, add2_i[28], n221);
  nand U304 ( n293, n295, n294);
  nand U305 ( n301, n303, n302);
  nand U306 ( n303, add2_i[10], n304);
  nand U307 ( n242, n244, n243);
  nand U308 ( n244, n245, add2_i[23]);
  or U309 ( n272, n273, add1_i[18]);
  nand U310 ( n264, n270, n269);
  nand U311 ( n261, add1_i[19], n264);
  nand U312 ( n231, add1_i[26], n338);
  nand U313 ( n246, n249, n248);
  nand U314 ( n273, n275, n274);
  nand U315 ( n274, add1_i[17], n277);
  nand U316 ( n204, add1_i[31], n333);
  nand U317 ( n208, add1_i[30], n337);
  nand U318 ( n253, add1_i[21], n256);
  nand U319 ( n277, n279, n278);
  nand U320 ( n207, n209, n208);
  nand U321 ( n211, n212, n213);
  nand U322 ( n234, n235, n236);
  nand U323 ( n256, n257, n258);
  nand U324 ( n281, n283, n282);
  nand U325 ( n282, n285, add1_i[15]);
  or U326 ( n305, n306, add1_i[10]);
  nand U327 ( n302, add1_i[10], n306);
  xnor U328 ( n188, n314, add1_i[8]);
  nand U329 ( n235, add1_i[25], n238);
  nand U330 ( n248, add1_i[22], n252);
  or U331 ( n251, n252, add1_i[22]);
  nand U332 ( n286, add1_i[14], n289);
  nand U333 ( n294, add1_i[12], n297);
  nand U334 ( n306, n308, n307);
  nand U335 ( n311, n312, n313, add1_i[8]);
  nand U336 ( n314, n313, n312);
  nor U337 ( result_o[6], n196, n357);
  xnor U338 ( result_o[27], add2_i[27], n230);
  not U339 ( n180, n357);
  nand U340 ( n219, add1_i[28], n227);
  or U341 ( n229, n230, n186);
  nand U342 ( n226, n231, n232);
  nand U343 ( n238, n239, n240);
  nand U344 ( n252, n254, n253);
  nand U345 ( n285, n287, n286);
  nand U346 ( n289, n291, n290);
  nand U347 ( n318, n181, n357);
  nand U348 ( n192, n319, n320);
  nand U349 ( result_o[32], n204, n205);
  nor U350 ( result_o[5], n332, n181);
  nand U351 ( n205, add2_i[31], n206);
  nor U352 ( n197, n332, n193);
  nor U353 ( n191, n193, n332, n180);
  nand U354 ( n227, n229, n225);
  nand U355 ( n222, n223, n224);
  nand U356 ( n224, n225, n186);
  nand U357 ( n243, add1_i[23], n246);
  or U358 ( n245, n246, add1_i[23]);
  nand U359 ( n258, add1_i[20], n259);
  nand U360 ( n257, add2_i[20], n260);
  nand U361 ( n259, n261, n262);
  nand U362 ( n278, add1_i[16], n281);
  nand U363 ( n283, add2_i[15], n284);
  nand U364 ( n297, n299, n298);
  nand U365 ( n310, n188, add2_i[8]);
  nor U366 ( result_o[2], n216, n353, n218);
  nand U367 ( n209, add2_i[30], n210);
  nand U368 ( n213, add2_i[29], n214);
  or U369 ( n223, n341, add1_i[27]);
  nand U370 ( n225, add1_i[27], n341);
  xnor U371 ( n230, n226, add1_i[27]);
  nand U372 ( n232, add2_i[26], n233);
  nand U373 ( n236, add2_i[25], n237);
  nand U374 ( n240, n241, add2_i[24]);
  nand U375 ( n254, n255, add2_i[21]);
  nand U376 ( n262, add2_i[19], n263);
  nand U377 ( n275, n276, add2_i[17]);
  nand U378 ( n279, n280, add2_i[16]);
  nand U379 ( n287, add2_i[14], n288);
  nand U380 ( n291, add2_i[13], n292);
  nand U381 ( n295, add2_i[12], n296);
  nand U382 ( n299, add2_i[11], n300);
  nand U383 ( n308, add2_i[9], n187);
endmodule
