// Verilog File 
module array_multiplier8_aor_enc128.bench (op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,product_o[0],product_o[1],product_o[2],product_o[3],product_o[4],
product_o[5],product_o[6],product_o[7],product_o[8],product_o[9],product_o[10],product_o[11],product_o[12],product_o[13],product_o[14],
product_o[15]);

input op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127;


output product_o[0], product_o[1], product_o[2], product_o[3], product_o[4], product_o[5], product_o[6], product_o[7], product_o[8], 
product_o[9], product_o[10], product_o[11], product_o[12], product_o[13], product_o[14], product_o[15];

wire xenc55, xenc35, n279, n280, xenc82, n281, xenc89, n284, n285, 
xenc47, xenc39, xenc6, xenc28, n296, n300, n318, xenc77, xenc95, xenc74, 
n319, n326, xenc4, n312, xenc106, n337, n353, n344, xenc38, xenc101, 
n350, n348, n378, n393, xenc68, n270, n397, n376, n351, xenc114, 
n370, n359, n371, n368, n405, xenc79, n374, xenc34, xenc20, n389, 
xenc41, n433, n430, xenc37, n417, n422, n411, n454, n410, xenc44, 
n416, xenc40, n453, n403, n401, n445, n473, xenc105, n437, xenc96, 
xenc69, n506, n507, n276, n508, n509, xenc9, n511, n474, n512, 
xenc86, n510, n514, n466, n452, xenc63, n463, xenc76, xenc25, n502, 
xenc93, xenc124, n540, n555, n556, n495, xenc110, xenc126, xenc85, n559, 
n527, n529, n580, xenc12, n592, n523, n530, n283, n255, n288, 
xenc56, n407, n408, n364, xenc30, n338, n521, xenc48, n259, n258, 
n267, n395, n396, n582, n583, n581, xenc119, xenc117, n383, n446, 
n404, n420, n423, n352, n325, n343, n341, xenc127, n517, xenc67, 
n442, n272, n443, xenc112, n441, xenc121, xenc13, xenc15, n363, n406, 
xenc122, n398, n356, n358, n306, n327, n311, xenc98, xenc11, n576, 
xenc64, n552, xenc53, n579, n584, n585, n541, n586, n587, n515, 
n460, n459, n457, xenc8, n503, n485, xenc1, n505, n390, n266, 
n391, n392, n588, xenc71, xenc87, n591, n589, n293, n301, n299, 
n292, xenc19, n332, xenc24, xenc27, n330, n360, n382, n261, n384, 
xenc26, n496, n480, n497, n498, n569, xenc21, n547, n571, n572, 
n570, n484, xenc97, n273, n486, xenc31, n551, xenc111, n277, n553, 
xenc54, xenc23, n438, n394, n439, n440, n548, n549, n550, n481, 
n482, n483, n488, n431, xenc116, n451, n537, xenc108, n539, n538, 
n399, n400, n402, n346, n347, n324, n349, n447, n448, xenc81, 
n450, n354, n355, n357, n427, xenc50, n429, n428, xenc60, n605, 
n499, n500, xenc103, n501, n477, n478, n479, n525, n526, n528, 
n386, xenc70, n263, xenc0, xenc88, xenc46, xenc49, n387, n388, xenc115, 
n373, n372, xenc75, n375, n566, xenc92, n543, xenc43, n567, n568, 
xenc109, xenc125, n432, n470, xenc52, n471, n472, n379, n380, n264, 
xenc72, n381, xenc65, n493, n475, n492, n494, n534, n535, n536, 
n320, n321, n317, xenc16, n322, n323, xenc62, xenc78, n465, n531, 
xenc73, n532, n533, n461, n462, n464, n313, n314, n298, xenc58, 
n316, n563, n564, n557, n565, xenc113, n425, n377, n424, n426, 
n339, xenc66, n342, n340, n418, xenc99, xenc51, n419, n421, n361, 
n362, n331, n328, xenc2, n305, n329, xenc104, xenc120, n303, n302, 
n333, xenc32, n336, n334, n412, n413, n365, n415, n366, n367, 
n369, n307, n308, n310, n560, n561, n562, n294, n295, n297, 
n289, n290, n287, n455, n456, n458, xenc57, xenc36, n519, n522, 
n520, xenc90, n603, n602, xenc5, n604, n593, xenc29, n595, n594, 
xenc94, n574, n573, n575, xenc107, xenc45, n489, n491, n490, xenc102, 
xenc59, n467, xenc18, n468, n469, n599, n600, n601, xenc14, xenc123, 
n434, xenc80, n435, n436, xenc33, n545, n504, n544, xenc42, n546, 
n596, n597, n598, xenc61, n409, xenc7, n345, xenc83, n265, xenc118, 
n262, xenc3, n577, xenc22, n516, n518, n256, n554, xenc17, n286, 
n578, xenc84, n487, n444, n524, n257, n269, n590, n449, n558, 
n513, n476, n414, n260, n542, n304, n268, n385, n606, xenc100, 
xenc91, n607, n335, n309, n271, xenc10, n291, n282, n608, n315;

xor g0(product_o[7], xenc55, xenc35);
xor g1(xenc82, n279, n280);
xor g2(product_o[1], n281, xenc89);
xor g3(product_o[14], n284, n285);
xor g4(xenc6, xenc47, xenc39);
xor g5(n300, xenc28, n296);
xor g6(product_o[12], n318, xenc77);
xor g7(n319, xenc95, xenc74);
xor g8(n318, n326, xenc4);
xor g9(n326, n312, xenc106);
xor g10(n344, n337, n353);
xor g11(product_o[10], xenc38, xenc101);
xor g12(n378, n350, n348);
xor g13(n270, n393, xenc68);
xor g14(n351, n397, n376);
xor g15(n359, xenc114, n370);
xor g16(n405, n371, n368);
xor g17(n397, xenc79, n374);
xor g18(n389, xenc34, xenc20);
xor g19(n430, xenc41, n433);
xor g20(n422, xenc37, n417);
xor g21(n417, n411, n454);
xor g22(n454, n410, xenc44);
xor g23(n453, n416, xenc40);
xor g24(n445, n403, n401);
xor g25(n437, n473, xenc105);
xor g26(n473, xenc96, xenc69);
xor g27(n276, n506, n507);
xor g28(n507, n508, n509);
xor g29(n474, xenc9, n511);
xor g30(n510, n512, xenc86);
xor g31(n452, n514, n466);
xor g32(n514, xenc63, n463);
xor g33(n502, xenc76, xenc25);
xor g34(n540, xenc93, xenc124);
xor g35(n495, n555, n556);
xor g36(n555, xenc110, xenc126);
xor g37(n511, xenc85, n559);
xor g38(n559, n527, n529);
xor g39(n280, n580, xenc12);
xor g40(n530, n592, n523);
not g41(n255, n283);
nor g42(n283, n288, xenc56);
nand g43(n364, n407, n408);
nand g44(n408, xenc44, n410);
nand g45(n407, xenc44, n411);
xnor g46(n353, xenc30, n338);
xnor g47(n592, n521, xenc48);
nor g48(n267, n259, n258, xenc35);
xnor g49(n393, n395, n396);
xnor g50(n581, n582, n583);
xnor g51(n383, xenc119, xenc117);
xnor g52(n404, n422, n446);
xnor g53(n446, n420, n423);
xnor g54(n325, n352, n344);
xnor g55(n352, n343, n341);
nor g56(n410, xenc127, n517);
xnor g57(n272, xenc67, n442);
xnor g58(n441, n443, xenc112);
xnor g59(n370, xenc121, xenc13);
xnor g60(n406, xenc15, n363);
xnor g61(n376, xenc122, n398);
xnor g62(n398, n356, n358);
xnor g63(n311, n306, n327);
xnor g64(n327, xenc98, xenc11);
xnor g65(n552, n576, xenc64);
xnor g66(n576, xenc53, n579);
xnor g67(n541, n584, n585);
xnor g68(n584, n586, n587);
xnor g69(n466, n515, n460);
xnor g70(n515, n459, n457);
xnor g71(n485, xenc8, n503);
xnor g72(n503, xenc1, n505);
xnor g73(n266, n389, n390);
xnor g74(n390, n391, n392);
xnor g75(n556, n588, xenc71);
xnor g76(n589, xenc87, n591);
xnor g77(n299, n293, n301);
xnor g78(n301, n292, xenc19);
xnor g79(n337, n332, xenc24);
xnor g80(n360, xenc27, n330);
xnor g81(n261, n382, n383);
xnor g82(n382, n384, xenc26);
xnor g83(n480, n495, n496);
xnor g84(n496, n497, n498);
xnor g85(n547, n569, xenc21);
xnor g86(n570, n571, n572);
xnor g87(n273, n484, xenc97);
xnor g88(n484, n486, xenc31);
xnor g89(n277, n551, xenc111);
xnor g90(n551, n553, xenc54);
xnor g91(n394, xenc23, n438);
xnor g92(n438, n439, n440);
xnor g93(n506, n547, n548);
xnor g94(n548, n549, n550);
xnor g95(n442, n480, n481);
xnor g96(n481, n482, n483);
xnor g97(n431, n452, n488);
xnor g98(n488, xenc116, n451);
nand g99(n498, n537, xenc108);
or g100(n537, n505, xenc1);
nand g101(n538, xenc8, n539);
nand g102(n539, xenc1, n505);
nand g103(n358, n399, n400);
nand g104(n399, xenc117, n403);
nand g105(n400, n401, n402);
or g106(n402, n403, xenc117);
nand g107(n324, n346, n347);
nand g108(n346, xenc38, n350);
nand g109(n347, n348, n349);
or g110(n349, n350, xenc38);
nand g111(n423, n447, n448);
nand g112(n447, n452, n451);
nand g113(n448, xenc116, xenc81);
or g114(n450, n451, n452);
nand g115(n338, n354, n355);
nand g116(n354, xenc122, n358);
nand g117(n355, n356, n357);
or g118(n357, n358, xenc122);
and g119(n384, n427, xenc50);
or g120(n427, n392, n391);
nand g121(n428, n389, n429);
nand g122(n429, n391, n392);
and g123(n579, xenc60, n583);
nand g124(n605, n582, n580);
and g125(n482, n499, n500);
or g126(n499, n486, xenc31);
nand g127(n500, xenc97, xenc103);
nand g128(n501, n486, xenc31);
and g129(n439, n477, n478);
or g130(n477, n443, xenc112);
nand g131(n478, n442, n479);
nand g132(n479, n443, xenc112);
and g133(n459, n525, n526);
or g134(n525, xenc85, n529);
nand g135(n526, n527, n528);
nand g136(n528, n529, xenc85);
and g137(n263, n386, xenc70);
nand g138(n386, xenc0, xenc88);
nand g139(n387, xenc46, xenc49);
or g140(n388, xenc0, xenc88);
and g141(n343, xenc115, n373);
nand g142(n372, n376, xenc79);
nand g143(n373, n374, xenc75);
or g144(n375, n376, xenc79);
nand g145(n543, n566, xenc92);
or g146(n566, n550, n549);
nand g147(n567, n547, xenc43);
nand g148(n568, n549, n550);
nor g149(product_o[15], n259, n283, xenc127);
nand g150(n432, xenc109, xenc125);
or g151(n470, n440, n439);
nand g152(n471, xenc23, xenc52);
nand g153(n472, n439, n440);
nand g154(n350, n379, n380);
or g155(n379, n264, xenc72);
nand g156(n380, n261, n381);
nand g157(n381, xenc72, n264);
nand g158(n475, xenc65, n493);
or g159(n492, n483, n482);
nand g160(n493, n480, n494);
nand g161(n494, n482, n483);
nand g162(n512, n534, n535);
nand g163(n534, n495, n498);
nand g164(n535, n497, n536);
or g165(n536, n498, n495);
nand g166(n317, n320, n321);
nand g167(n320, xenc16, n324);
nand g168(n321, n322, n323);
or g169(n323, n324, xenc16);
nand g170(n465, xenc62, xenc78);
nand g171(n531, n511, n512);
nand g172(n532, xenc86, xenc73);
or g173(n533, n512, n511);
nand g174(n416, n461, n462);
nand g175(n461, n466, xenc63);
nand g176(n462, n463, n464);
or g177(n464, xenc63, n466);
nand g178(n298, n313, n314);
nand g179(n313, n318, xenc95);
nand g180(n314, xenc74, xenc58);
or g181(n316, xenc95, n318);
nand g182(n557, n563, n564);
nand g183(n563, xenc25, xenc124);
nand g184(n564, xenc93, n565);
or g185(n565, xenc124, xenc25);
nand g186(n377, xenc113, n425);
or g187(n424, n383, n384);
nand g188(n425, xenc26, n426);
nand g189(n426, n383, n384);
nand g190(n312, n339, xenc66);
or g191(n339, n344, n343);
nand g192(n340, n341, n342);
nand g193(n342, n343, n344);
nand g194(n371, n418, xenc99);
nand g195(n418, n422, n423);
nand g196(n419, n420, xenc51);
or g197(n421, n422, n423);
nand g198(n331, n361, n362);
nand g199(n362, n363, xenc15);
nand g200(n361, n363, xenc121);
nand g201(n305, n328, xenc2);
nand g202(n329, n330, xenc27);
nand g203(n328, n330, n332);
nand g204(n292, xenc104, xenc120);
nand g205(n303, xenc11, xenc98);
nand g206(n302, xenc11, n306);
nand g207(n306, n333, xenc32);
nand g208(n333, n337, n338);
nand g209(n334, xenc30, n336);
or g210(n336, n337, n338);
nand g211(n365, n412, n413);
nand g212(n412, n417, n416);
nand g213(n413, xenc40, n415);
or g214(n415, n416, n417);
nand g215(n332, n366, n367);
nand g216(n366, n370, n371);
nand g217(n367, n368, n369);
or g218(n369, n370, n371);
nand g219(n293, n307, n308);
nand g220(n307, xenc4, n312);
nand g221(n308, xenc106, n310);
or g222(n310, xenc4, n312);
and g223(n529, n560, n561);
nand g224(n560, n556, xenc110);
nand g225(n561, xenc126, n562);
or g226(n562, xenc110, n556);
nand g227(n288, n294, n295);
nand g228(n294, xenc39, xenc28);
nand g229(n295, n296, n297);
or g230(n297, xenc28, xenc39);
nand g231(n583, product_o[0], n580);
nand g232(n287, n289, n290);
nand g233(n290, xenc19, n292);
nand g234(n289, xenc19, n293);
nand g235(n411, n455, n456);
or g236(n455, n460, n459);
nand g237(n456, n457, n458);
nand g238(n458, n459, n460);
and g239(n517, xenc57, xenc36);
nand g240(n519, xenc48, n523);
nand g241(n520, n521, n522);
or g242(n522, n523, xenc48);
and g243(n569, xenc90, n603);
or g244(n602, xenc64, n579);
nand g245(n603, xenc53, xenc5);
nand g246(n604, n579, xenc64);
nand g247(n523, n593, xenc29);
or g248(n593, n591, n588);
nand g249(n594, xenc87, n595);
nand g250(n595, n588, n591);
and g251(n549, xenc94, n574);
or g252(n573, n553, xenc54);
nand g253(n574, xenc111, n575);
nand g254(n575, n553, xenc54);
nand g255(n451, xenc107, xenc45);
nand g256(n489, xenc105, xenc96);
nand g257(n490, xenc69, n491);
or g258(n491, xenc96, xenc105);
nand g259(n403, xenc102, xenc59);
nand g260(n467, xenc20, xenc41);
nand g261(n468, n433, xenc18);
or g262(n469, xenc41, xenc20);
nand g263(n585, n599, n600);
or g264(n599, n572, n569);
nand g265(n600, n571, n601);
nand g266(n601, n569, n572);
and g267(n391, xenc14, xenc123);
or g268(n434, n395, n396);
nand g269(n435, xenc68, xenc80);
nand g270(n436, n395, n396);
and g271(n504, xenc33, n545);
or g272(n544, n508, n509);
nand g273(n545, n506, xenc42);
nand g274(n546, n508, n509);
and g275(n588, n596, n597);
nand g276(n596, n586, n585);
nand g277(n597, n587, n598);
or g278(n598, n585, n586);
nor g279(n409, xenc127, xenc61);
xnor g280(product_o[11], xenc16, xenc7);
xnor g281(n345, n322, n324);
xnor g282(product_o[8], xenc83, xenc46);
xnor g283(n265, xenc0, xenc88);
xnor g284(product_o[9], n261, xenc118);
xnor g285(n262, xenc72, n264);
nor g286(n279, xenc61, n258);
nand g287(n553, op2_i[2], n280, op1_i[0]);
nand g288(n486, op1_i[0], n276, op2_i[4]);
nand g289(n395, op1_i[0], xenc3, op2_i[6]);
nand g290(n443, op2_i[5], op1_i[0], n273);
nand g291(n577, op1_i[2], op2_i[1]);
nand g292(n572, op2_i[1], op1_i[3]);
nand g293(n550, op1_i[2], op2_i[2]);
nand g294(n460, xenc22, n516);
nand g295(n516, n517, n518);
not g296(n256, n410);
nand g297(n518, op1_i[7], op2_i[1]);
nand g298(n554, op1_i[1], op2_i[2]);
nand g299(n508, op2_i[3], op1_i[0], n277);
and g300(n580, op2_i[1], op1_i[1]);
and g301(n586, op2_i[1], op1_i[4]);
and g302(n587, op2_i[0], op1_i[5]);
nand g303(n285, op2_i[7], op1_i[7]);
nand g304(n284, n255, xenc17);
nand g305(n286, xenc56, n288);
and g306(n582, op2_i[0], op1_i[2]);
and g307(n578, op2_i[0], op1_i[3]);
and g308(n571, op2_i[0], op1_i[4]);
and g309(xenc84, op1_i[0], op2_i[0]);
nand g310(n505, op2_i[3], op1_i[2]);
nand g311(n591, op2_i[1], op1_i[5]);
nand g312(n483, op2_i[4], op1_i[2]);
nand g313(n440, op2_i[5], op1_i[2]);
nand g314(n487, op2_i[4], op1_i[1]);
nand g315(n444, op2_i[5], op1_i[1]);
and g316(n524, op2_i[1], op1_i[6]);
not g317(n257, op1_i[7]);
nand g318(n509, op2_i[3], op1_i[1]);
and g319(n457, op2_i[2], op1_i[6]);
nand g320(n269, op2_i[7], op1_i[0]);
and g321(n590, op2_i[0], op1_i[6]);
and g322(n497, op2_i[3], op1_i[3]);
and g323(n521, op1_i[7], op2_i[0]);
and g324(n449, op2_i[4], op1_i[4]);
and g325(n558, op1_i[4], op2_i[2]);
and g326(n513, op2_i[3], op1_i[4]);
and g327(n476, op2_i[4], op1_i[3]);
and g328(n463, op2_i[3], op1_i[5]);
and g329(n414, op2_i[3], op1_i[6]);
not g330(n260, op2_i[2]);
and g331(n542, op1_i[3], op2_i[2]);
and g332(n527, op1_i[5], op2_i[2]);
nand g333(n392, op2_i[6], op1_i[2]);
nand g334(n264, op2_i[7], op1_i[2]);
and g335(n363, op2_i[3], op1_i[7]);
and g336(n330, op2_i[4], op1_i[7]);
and g337(n304, op2_i[5], op1_i[7]);
nand g338(n396, op2_i[6], op1_i[1]);
and g339(n268, op2_i[7], op1_i[1]);
and g340(n385, op2_i[6], op1_i[3]);
and g341(n341, op2_i[6], op1_i[5]);
xnor g342(xenc100, n606, n276);
nand g343(n606, op1_i[0], op2_i[4]);
xnor g344(product_o[5], n273, xenc91);
nand g345(n607, op1_i[0], op2_i[5]);
and g346(n420, op2_i[4], op1_i[5]);
and g347(n356, op2_i[5], op1_i[5]);
and g348(n335, op2_i[5], op1_i[6]);
and g349(n322, op2_i[7], op1_i[4]);
not g350(n259, op2_i[7]);
and g351(n433, op2_i[5], op1_i[3]);
and g352(n401, op2_i[5], op1_i[4]);
and g353(n368, op2_i[4], op1_i[6]);
and g354(n374, op2_i[6], op1_i[4]);
and g355(n348, op2_i[7], op1_i[3]);
and g356(n309, op2_i[6], op1_i[6]);
not g357(n258, op1_i[0]);
xnor g358(xenc10, n271, xenc3);
nand g359(n271, op2_i[6], op1_i[0]);
and g360(n291, op2_i[6], op1_i[7]);
nand g361(n281, op2_i[0], op1_i[1]);
nand g362(n282, op1_i[0], op2_i[1]);
xnor g363(product_o[3], n277, n608);
nand g364(n608, op1_i[0], op2_i[3]);
and g365(n315, op2_i[7], op1_i[5]);
and g366(n296, op2_i[7], op1_i[6]);
or g367(xenc0, n267, keyinput0);
and g368(xenc1, n504, keyinput1);
and g369(xenc2, n329, keyinput2);
and g370(xenc3, n272, keyinput3);
or g371(xenc4, n311, keyinput4);
and g372(xenc5, n604, keyinput5);
or g373(product_o[13], xenc6, keyinput6);
or g374(xenc7, n345, keyinput7);
or g375(xenc8, n502, keyinput8);
or g376(xenc9, n510, keyinput9);
and g377(product_o[6], xenc10, keyinput10);
or g378(xenc11, n304, keyinput11);
or g379(xenc12, n581, keyinput12);
or g380(xenc13, n406, keyinput13);
or g381(xenc14, n434, keyinput14);
or g382(xenc15, n364, keyinput15);
or g383(xenc16, n325, keyinput16);
and g384(xenc17, n286, keyinput17);
and g385(xenc18, n469, keyinput18);
or g386(xenc19, n291, keyinput19);
and g387(xenc20, n431, keyinput20);
and g388(xenc21, n570, keyinput21);
or g389(xenc22, n256, keyinput22);
or g390(xenc23, n437, keyinput23);
and g391(xenc24, n360, keyinput24);
or g392(xenc25, n541, keyinput25);
or g393(xenc26, n385, keyinput26);
and g394(xenc27, n331, keyinput27);
and g395(xenc28, n298, keyinput28);
or g396(xenc29, n594, keyinput29);
or g397(xenc30, n335, keyinput30);
or g398(xenc31, n487, keyinput31);
or g399(xenc32, n334, keyinput32);
or g400(xenc33, n544, keyinput33);
and g401(xenc34, n430, keyinput34);
and g402(xenc35, n270, keyinput35);
or g403(xenc36, n520, keyinput36);
or g404(xenc37, n453, keyinput37);
and g405(xenc38, n351, keyinput38);
and g406(xenc39, n299, keyinput39);
and g407(xenc40, n414, keyinput40);
and g408(xenc41, n432, keyinput41);
and g409(xenc42, n546, keyinput42);
and g410(xenc43, n568, keyinput43);
or g411(xenc44, n409, keyinput44);
or g412(xenc45, n490, keyinput45);
or g413(xenc46, n266, keyinput46);
and g414(xenc47, n300, keyinput47);
or g415(xenc48, n524, keyinput48);
or g416(xenc49, n388, keyinput49);
or g417(xenc50, n428, keyinput50);
or g418(xenc51, n421, keyinput51);
and g419(xenc52, n472, keyinput52);
and g420(xenc53, n578, keyinput53);
or g421(xenc54, n554, keyinput54);
and g422(xenc55, n269, keyinput55);
and g423(xenc56, n287, keyinput56);
and g424(xenc57, n519, keyinput57);
or g425(xenc58, n316, keyinput58);
and g426(xenc59, n468, keyinput59);
or g427(xenc60, n605, keyinput60);
and g428(xenc61, n260, keyinput61);
or g429(xenc62, n531, keyinput62);
and g430(xenc63, n465, keyinput63);
or g431(xenc64, n577, keyinput64);
or g432(xenc65, n492, keyinput65);
and g433(xenc66, n340, keyinput66);
and g434(xenc67, n441, keyinput67);
and g435(xenc68, n394, keyinput68);
and g436(xenc69, n476, keyinput69);
and g437(xenc70, n387, keyinput70);
or g438(xenc71, n589, keyinput71);
and g439(xenc72, n263, keyinput72);
and g440(xenc73, n533, keyinput73);
or g441(xenc74, n315, keyinput74);
or g442(xenc75, n375, keyinput75);
and g443(xenc76, n540, keyinput76);
and g444(xenc77, n319, keyinput77);
or g445(xenc78, n532, keyinput78);
or g446(xenc79, n377, keyinput79);
and g447(xenc80, n436, keyinput80);
and g448(xenc81, n450, keyinput81);
or g449(product_o[2], xenc82, keyinput82);
and g450(xenc83, n265, keyinput83);
or g451(product_o[0], xenc84, keyinput84);
and g452(xenc85, n530, keyinput85);
and g453(xenc86, n513, keyinput86);
or g454(xenc87, n590, keyinput87);
and g455(xenc88, n268, keyinput88);
or g456(xenc89, n282, keyinput89);
or g457(xenc90, n602, keyinput90);
or g458(xenc91, n607, keyinput91);
or g459(xenc92, n567, keyinput92);
and g460(xenc93, n542, keyinput93);
or g461(xenc94, n573, keyinput94);
and g462(xenc95, n317, keyinput95);
and g463(xenc96, n475, keyinput96);
or g464(xenc97, n485, keyinput97);
and g465(xenc98, n305, keyinput98);
and g466(xenc99, n419, keyinput99);
and g467(product_o[4], xenc100, keyinput100);
or g468(xenc101, n378, keyinput101);
or g469(xenc102, n467, keyinput102);
and g470(xenc103, n501, keyinput103);
or g471(xenc104, n302, keyinput104);
and g472(xenc105, n474, keyinput105);
and g473(xenc106, n309, keyinput106);
or g474(xenc107, n489, keyinput107);
or g475(xenc108, n538, keyinput108);
or g476(xenc109, n470, keyinput109);
or g477(xenc110, n557, keyinput110);
or g478(xenc111, n552, keyinput111);
and g479(xenc112, n444, keyinput112);
and g480(xenc113, n424, keyinput113);
or g481(xenc114, n405, keyinput114);
or g482(xenc115, n372, keyinput115);
and g483(xenc116, n449, keyinput116);
or g484(xenc117, n404, keyinput117);
and g485(xenc118, n262, keyinput118);
and g486(xenc119, n445, keyinput119);
or g487(xenc120, n303, keyinput120);
or g488(xenc121, n365, keyinput121);
or g489(xenc122, n359, keyinput122);
and g490(xenc123, n435, keyinput123);
or g491(xenc124, n543, keyinput124);
and g492(xenc125, n471, keyinput125);
or g493(xenc126, n558, keyinput126);
or g494(xenc127, n257, keyinput127);
endmodule
