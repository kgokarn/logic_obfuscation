module carry_lookahead_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136;

  xor U126 ( result_o[9], n61, n62);
  xor U127 ( n62, add2_i[9], add1_i[9]);
  xor U128 ( result_o[8], n63, n64);
  xor U129 ( n64, add2_i[8], add1_i[8]);
  xor U130 ( result_o[7], n65, n66);
  xor U131 ( n66, add2_i[7], add1_i[7]);
  xor U132 ( result_o[6], n67, n68);
  xor U133 ( n68, add2_i[6], add1_i[6]);
  xor U134 ( result_o[5], n69, n70);
  xor U135 ( n70, add2_i[5], add1_i[5]);
  xor U136 ( result_o[4], n71, n72);
  xor U137 ( n72, add2_i[4], add1_i[4]);
  xor U138 ( result_o[3], n73, n74);
  xor U139 ( n74, add2_i[3], add1_i[3]);
  xor U140 ( result_o[2], n75, n76);
  xor U141 ( n76, add2_i[2], add1_i[2]);
  xor U142 ( result_o[1], n77, n78);
  xor U143 ( n78, add2_i[1], add1_i[1]);
  xor U144 ( result_o[15], n82, n83);
  xor U145 ( n83, add2_i[15], add1_i[15]);
  xor U146 ( result_o[14], n87, n88);
  xor U147 ( n88, add2_i[14], add1_i[14]);
  xor U148 ( result_o[13], n92, n93);
  xor U149 ( n93, add2_i[13], add1_i[13]);
  xor U150 ( result_o[12], n97, n98);
  xor U151 ( n98, add2_i[12], add1_i[12]);
  xor U152 ( result_o[11], n102, n103);
  xor U153 ( n103, add2_i[11], add1_i[11]);
  xor U154 ( result_o[10], n107, n108);
  xor U155 ( n108, add2_i[10], add1_i[10]);
  or U156 ( n77, add2_i[0], add1_i[0]);
  nand U157 ( n75, n133, n134);
  nand U158 ( n133, add1_i[1], n77);
  nand U159 ( n134, add2_i[1], n135);
  or U160 ( n135, n77, add1_i[1]);
  nand U161 ( n73, n130, n131);
  nand U162 ( n130, add1_i[2], n75);
  nand U163 ( n131, add2_i[2], n132);
  or U164 ( n132, n75, add1_i[2]);
  nand U165 ( n92, n94, n95);
  nand U166 ( n94, add1_i[12], n97);
  nand U167 ( n95, add2_i[12], n96);
  or U168 ( n96, n97, add1_i[12]);
  nand U169 ( n87, n89, n90);
  nand U170 ( n89, add1_i[13], n92);
  nand U171 ( n90, add2_i[13], n91);
  or U172 ( n91, n92, add1_i[13]);
  nand U173 ( n82, n84, n85);
  nand U174 ( n84, add1_i[14], n87);
  nand U175 ( n85, add2_i[14], n86);
  or U176 ( n86, n87, add1_i[14]);
  nand U177 ( n71, n127, n128);
  nand U178 ( n127, add1_i[3], n73);
  nand U179 ( n128, add2_i[3], n129);
  or U180 ( n129, n73, add1_i[3]);
  nand U181 ( n69, n124, n125);
  nand U182 ( n124, add1_i[4], n71);
  nand U183 ( n125, add2_i[4], n126);
  or U184 ( n126, n71, add1_i[4]);
  nand U185 ( n67, n121, n122);
  nand U186 ( n121, add1_i[5], n69);
  nand U187 ( n122, add2_i[5], n123);
  or U188 ( n123, n69, add1_i[5]);
  nand U189 ( n65, n118, n119);
  nand U190 ( n118, add1_i[6], n67);
  nand U191 ( n119, add2_i[6], n120);
  or U192 ( n120, n67, add1_i[6]);
  nand U193 ( n63, n115, n116);
  nand U194 ( n115, add1_i[7], n65);
  nand U195 ( n116, add2_i[7], n117);
  or U196 ( n117, n65, add1_i[7]);
  nand U197 ( n61, n112, n113);
  nand U198 ( n112, add1_i[8], n63);
  nand U199 ( n113, add2_i[8], n114);
  or U200 ( n114, n63, add1_i[8]);
  nand U201 ( n107, n109, n110);
  nand U202 ( n109, add1_i[9], n61);
  nand U203 ( n110, add2_i[9], n111);
  or U204 ( n111, n61, add1_i[9]);
  nand U205 ( n102, n104, n105);
  nand U206 ( n104, add1_i[10], n107);
  nand U207 ( n105, add2_i[10], n106);
  or U208 ( n106, n107, add1_i[10]);
  nand U209 ( n97, n99, n100);
  nand U210 ( n99, add1_i[11], n102);
  nand U211 ( n100, add2_i[11], n101);
  or U212 ( n101, n102, add1_i[11]);
  nand U213 ( result_o[16], n79, n80);
  nand U214 ( n79, add1_i[15], n82);
  nand U215 ( n80, add2_i[15], n81);
  or U216 ( n81, n82, add1_i[15]);
  nand U217 ( result_o[0], n77, n136);
  nand U218 ( n136, add2_i[0], add1_i[0]);
endmodule
