library verilog;
use verilog.vl_types.all;
entity almost_correct_adder16_tb is
end almost_correct_adder16_tb;
