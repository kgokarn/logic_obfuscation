// Verilog File 
module broken_array_multiplier8_xor_enc128.bench (op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,product_o[0],product_o[1],product_o[2],product_o[3],product_o[4],
product_o[5],product_o[6],product_o[7],product_o[8],product_o[9],product_o[10],product_o[11],product_o[12],product_o[13],product_o[14],
product_o[15]);

input op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127;


output product_o[0], product_o[1], product_o[2], product_o[3], product_o[4], product_o[5], product_o[6], product_o[7], product_o[8], 
product_o[9], product_o[10], product_o[11], product_o[12], product_o[13], product_o[14], product_o[15];

wire n203, n204, xenc0, xenc111, n222, n223, xenc12, xenc21, n230, 
xenc18, n237, n229, n231, n239, n236, xenc97, n238, n258, xenc64, 
xenc88, n256, xenc58, xenc109, xenc125, xenc30, xenc1, n279, n283, xenc50, 
n298, n275, n325, xenc68, n208, xenc7, n328, n347, n348, n330, 
xenc84, n350, n355, xenc105, n319, xenc16, n312, n296, xenc34, n361, 
n307, n313, n310, n359, xenc28, xenc51, xenc75, n386, n383, xenc107, 
xenc22, n352, n392, n393, n390, xenc89, xenc92, n341, n402, n373, 
xenc11, xenc86, xenc70, n442, n384, n443, n444, xenc31, n445, n398, 
n406, n408, n461, xenc103, n429, n467, n468, n465, xenc10, xenc3, 
n409, xenc8, xenc6, n219, n221, n357, xenc118, n356, n400, xenc99, 
n399, xenc63, n464, n462, xenc14, n265, n276, n273, n297, n333, 
n289, n293, xenc80, xenc78, xenc46, n441, n455, n456, n436, n457, 
n458, n250, xenc48, n257, xenc26, n251, n259, n290, n282, xenc96, 
n264, n334, n335, n295, n320, n321, n336, n291, xenc94, n294, 
n292, xenc67, xenc71, n260, n263, n261, xenc87, n420, n372, n419, 
n421, n284, xenc120, n281, xenc55, n288, xenc113, n287, n285, n277, 
xenc121, xenc53, n278, n280, n252, n253, n255, xenc43, n375, n374, 
n376, xenc29, n450, n430, n449, xenc85, n451, n377, n378, n358, 
n342, n343, n379, n246, xenc20, xenc69, n247, n249, xenc77, xenc62, 
n225, n232, n235, n233, n452, n453, xenc36, xenc91, n454, n422, 
n423, n401, n424, n473, n474, xenc54, n475, xenc81, xenc49, n476, 
xenc110, n477, n478, n308, xenc40, xenc19, n309, n311, xenc27, n447, 
n446, n448, n302, xenc65, xenc106, xenc57, xenc108, xenc127, n469, n244, 
n266, n242, n245, n351, n214, xenc73, n354, xenc37, n212, n331, 
xenc60, n329, n394, n395, n216, xenc104, n397, xenc17, n435, n367, 
n403, n364, n366, n318, n340, n326, n428, n391, xenc23, xenc44, 
n360, xenc4, xenc116, n315, xenc9, n316, n317, xenc24, n405, n404, 
n407, xenc33, xenc38, n380, xenc32, n381, n382, xenc41, xenc90, n337, 
xenc102, n338, n339, xenc25, xenc123, n306, n368, n371, n369, n271, 
n272, n274, xenc119, n388, n349, n387, n389, n344, xenc15, n327, 
n346, n345, n322, n323, n205, n209, xenc82, xenc72, xenc45, n324, 
n300, n270, n432, xenc13, xenc47, n433, n434, xenc2, n268, n470, 
n471, n417, n472, xenc56, n314, xenc126, xenc112, n240, xenc93, n241, 
n243, xenc5, n227, n224, n226, n228, n425, n426, n385, xenc59, 
n427, n362, n363, n301, n365, n413, xenc114, n412, xenc66, n414, 
n416, n303, xenc52, n269, xenc124, n304, n305, xenc101, n207, xenc115, 
xenc35, n460, n481, n482, n479, n480, xenc83, n220, n485, xenc39, 
n466, n486, n459, n440, xenc74, n484, n483, n439, xenc79, n218, 
xenc117, n353, n437, xenc122, n396, n418, n438, n410, n202, n411, 
n431, n463, n415, xenc100, n267, n210, n332, n299, n206, n286, 
n262, n248, xenc42, n213, xenc95, n211, n370, n215, xenc61, n487, 
n254, n234, xenc76, xenc98;

xor g0(product_o[9], n203, n204);
xor g1(n203, xenc0, xenc111);
xor g2(product_o[14], n222, n223);
xor g3(product_o[13], xenc12, xenc21);
xor g4(n237, n230, xenc18);
xor g5(n239, n229, n231);
xor g6(n238, n236, xenc97);
xor g7(xenc88, n258, xenc64);
xor g8(n258, n256, xenc58);
xor g9(xenc30, xenc109, xenc125);
xor g10(n283, xenc1, n279);
xor g11(n275, xenc50, n298);
xor g12(n208, n325, xenc68);
xor g13(n325, xenc7, n328);
xor g14(n330, n347, n348);
xor g15(n347, xenc84, n350);
xor g16(n319, n355, xenc105);
xor g17(n296, xenc16, n312);
xor g18(n307, xenc34, n361);
xor g19(n359, n313, n310);
xor g20(n348, xenc28, xenc51);
xor g21(n383, xenc75, n386);
xor g22(n352, xenc107, xenc22);
xor g23(n390, n392, n393);
xor g24(n341, xenc89, xenc92);
xor g25(n355, n402, n373);
xor g26(n402, xenc11, xenc86);
xor g27(n384, xenc70, n442);
xor g28(n442, n443, n444);
xor g29(n398, xenc31, n445);
xor g30(n445, n406, n408);
xor g31(n429, n461, xenc103);
xor g32(n465, n467, n468);
xor g33(n409, xenc10, xenc3);
nand g34(n219, xenc8, xenc6);
or g35(n221, xenc6, xenc8);
xnor g36(n356, n357, xenc118);
xnor g37(n399, n400, xenc99);
xnor g38(n462, xenc63, n464);
xnor g39(n265, xenc14, n275);
xnor g40(n297, n276, n273);
xnor g41(n289, n296, n333);
xnor g42(n333, n293, xenc80);
xnor g43(n441, xenc78, xenc46);
xnor g44(n436, n455, n456);
xnor g45(n455, n457, n458);
xnor g46(n257, n250, xenc48);
xnor g47(n259, xenc26, n251);
xnor g48(n282, n265, n290);
xnor g49(n290, xenc96, n264);
nand g50(n295, n334, n335);
or g51(n334, n319, n320);
nand g52(n335, n321, n336);
nand g53(n336, n320, n319);
nand g54(n264, n291, xenc94);
nand g55(n291, n296, xenc80);
nand g56(n292, n293, n294);
or g57(n294, xenc80, n296);
nand g58(n251, xenc67, xenc71);
nand g59(n260, n265, n264);
nand g60(n261, xenc96, n263);
or g61(n263, n264, n265);
nand g62(n372, xenc87, n420);
nand g63(n419, xenc89, xenc99);
nand g64(n420, n400, n421);
or g65(n421, xenc99, xenc89);
nand g66(n281, n284, xenc120);
nand g67(n284, xenc55, n288);
nand g68(n285, xenc113, n287);
or g69(n287, n288, xenc55);
nand g70(n256, n277, xenc121);
nand g71(n277, xenc109, xenc1);
nand g72(n278, n279, xenc53);
or g73(n280, xenc1, xenc109);
nand g74(n236, n252, n253);
nand g75(n252, xenc64, n256);
nand g76(n253, xenc58, n255);
or g77(n255, n256, xenc64);
nand g78(n313, xenc43, n375);
nand g79(n374, n355, xenc118);
nand g80(n375, n357, n376);
or g81(n376, n355, xenc118);
and g82(n444, xenc29, n450);
or g83(n449, n429, n430);
nand g84(n450, xenc85, n451);
nand g85(n451, n430, n429);
nand g86(n358, n377, n378);
or g87(n377, n341, n342);
nand g88(n378, n343, n379);
nand g89(n379, n342, n341);
and g90(n230, n246, xenc20);
nand g91(n246, n250, n251);
nand g92(n247, xenc26, xenc69);
or g93(n249, n250, n251);
nand g94(n225, xenc77, xenc62);
nand g95(n232, xenc21, n236);
nand g96(n233, xenc97, n235);
or g97(n235, n236, xenc21);
and g98(n430, n452, n453);
or g99(n452, xenc36, xenc91);
nand g100(n453, n436, n454);
nand g101(n454, xenc36, xenc91);
nand g102(n401, n422, n423);
nand g103(n422, xenc51, xenc75);
nand g104(n423, n386, n424);
or g105(n424, xenc75, xenc51);
nand g106(n468, n473, n474);
nand g107(n473, n461, n464);
nand g108(n474, xenc63, xenc54);
or g109(n475, n464, n461);
nand g110(n464, xenc81, xenc49);
nand g111(n476, n457, n456);
nand g112(n477, n458, xenc110);
or g113(n478, n456, n457);
and g114(n276, n308, xenc40);
nand g115(n308, n312, n313);
nand g116(n309, n310, xenc19);
or g117(n311, n312, n313);
and g118(n408, xenc27, n447);
or g119(n446, xenc70, n444);
nand g120(n447, n443, n448);
nand g121(n448, n444, xenc70);
xnor g122(n361, n302, xenc65);
xnor g123(n298, xenc106, xenc57);
xnor g124(n469, xenc108, xenc127);
xnor g125(n250, n244, n266);
xnor g126(n266, n242, n245);
xnor g127(n214, n351, n352);
xnor g128(n351, xenc73, n354);
xnor g129(n212, xenc37, n330);
xnor g130(n329, n331, xenc60);
xnor g131(n216, n394, n395);
xnor g132(n394, xenc104, n397);
xnor g133(n395, xenc17, n436);
xnor g134(n435, xenc36, xenc91);
xnor g135(n373, n367, n403);
xnor g136(n403, n364, n366);
xnor g137(n204, n318, n319);
xnor g138(n318, n320, n321);
xnor g139(n326, n340, n341);
xnor g140(n340, n342, n343);
xnor g141(n391, n428, n429);
xnor g142(n428, n430, xenc85);
xnor g143(n312, xenc23, n307);
xnor g144(n360, xenc44, xenc106);
nand g145(n288, xenc4, xenc116);
nand g146(n315, xenc111, xenc0);
nand g147(n316, n204, xenc9);
or g148(n317, xenc0, xenc111);
nand g149(n366, xenc24, n405);
or g150(n404, xenc31, n408);
nand g151(n405, n406, n407);
nand g152(n407, n408, xenc31);
and g153(n342, xenc33, xenc38);
nand g154(n380, n350, xenc84);
nand g155(n381, n348, xenc32);
or g156(n382, xenc84, n350);
and g157(n320, xenc41, xenc90);
nand g158(n337, n328, xenc7);
nand g159(n338, xenc68, xenc102);
or g160(n339, xenc7, n328);
and g161(n306, xenc25, xenc123);
nand g162(n368, n373, xenc11);
nand g163(n369, xenc86, n371);
or g164(n371, xenc11, n373);
and g165(n244, n271, n272);
or g166(n271, n275, n276);
nand g167(n272, n273, n274);
nand g168(n274, n275, n276);
nand g169(n349, xenc119, n388);
or g170(n387, xenc73, n354);
nand g171(n388, n352, n389);
nand g172(n389, xenc73, n354);
nand g173(n327, n344, xenc15);
nand g174(n344, n331, xenc60);
nand g175(n345, n330, n346);
or g176(n346, n331, xenc60);
nand g177(n205, n322, n323);
or g178(n322, n209, xenc82);
nand g179(n323, xenc72, xenc45);
nand g180(n324, n209, xenc82);
nand g181(n270, xenc65, n300);
nand g182(n300, xenc34, n302);
nand g183(n392, n432, xenc13);
or g184(n432, xenc104, n397);
nand g185(n433, n395, xenc47);
nand g186(n434, xenc104, n397);
and g187(n242, xenc106, xenc2);
nand g188(n268, xenc50, xenc57);
and g189(n417, n470, n471);
nand g190(n470, xenc46, n468);
nand g191(n471, n467, n472);
or g192(n472, n468, xenc46);
xnor g193(product_o[10], xenc55, xenc56);
xnor g194(n314, xenc113, n288);
nand g195(n229, xenc126, xenc112);
or g196(n240, n245, n244);
nand g197(n241, n242, xenc93);
nand g198(n243, n244, n245);
nand g199(n224, xenc5, n227);
or g200(n226, n231, n230);
nand g201(n227, n228, n229);
nand g202(n228, n230, n231);
nand g203(n385, n425, n426);
nand g204(n425, n393, n392);
nand g205(n426, xenc22, xenc59);
or g206(n427, n392, n393);
and g207(n301, n362, n363);
nand g208(n362, n367, n366);
nand g209(n363, n364, n365);
or g210(n365, n366, n367);
nand g211(n412, n413, xenc114);
or g212(n413, xenc127, xenc10);
nand g213(n414, xenc108, xenc66);
nand g214(n416, xenc10, xenc127);
and g215(n269, n303, xenc52);
or g216(n303, n307, xenc44);
nand g217(n304, xenc106, xenc124);
nand g218(n305, xenc44, n307);
xnor g219(product_o[8], xenc101, xenc72);
xnor g220(n207, n209, xenc82);
nand g221(n223, op2_i[7], op1_i[7]);
nand g222(n222, xenc115, xenc35);
and g223(n457, op2_i[2], n460, op1_i[2]);
xnor g224(n460, n481, n482);
nand g225(n481, op1_i[3], op2_i[1]);
and g226(n482, op1_i[4], op2_i[0]);
xnor g227(n456, n479, n480);
nand g228(n479, op1_i[4], op2_i[1]);
and g229(n480, op1_i[5], op2_i[0]);
nand g230(product_o[15], xenc35, xenc83);
nand g231(n220, op1_i[7], xenc115, op2_i[7]);
xnor g232(n466, n485, xenc39);
nand g233(n485, op1_i[6], op2_i[1]);
and g234(n486, op1_i[7], op2_i[0]);
xnor g235(n440, n459, n460);
nand g236(n459, op1_i[2], op2_i[2]);
xnor g237(n461, xenc74, n484);
nand g238(n483, op1_i[5], op2_i[1]);
and g239(n484, op1_i[6], op2_i[0]);
xnor g240(n218, n439, xenc79);
nand g241(n439, op1_i[1], op2_i[3]);
nand g242(n209, op1_i[0], xenc117, op2_i[7]);
nand g243(n353, op1_i[0], n216, op2_i[5]);
nand g244(n437, op2_i[3], xenc79, op1_i[1]);
nand g245(n396, op2_i[4], xenc122, op1_i[0]);
nand g246(n418, op2_i[2], op1_i[6]);
nand g247(n438, op2_i[3], op1_i[2]);
nand g248(n397, op2_i[4], op1_i[1]);
nand g249(n354, op2_i[5], op1_i[1]);
nand g250(n302, op1_i[7], n412);
and g251(n367, n302, n410);
nand g252(n410, n202, n411);
nand g253(n411, op2_i[2], op1_i[7]);
not g254(n202, n412);
and g255(n458, op1_i[3], op2_i[2]);
and g256(n431, op2_i[3], op1_i[3]);
and g257(n393, op2_i[4], op1_i[2]);
and g258(n350, op2_i[5], op1_i[2]);
and g259(n463, op1_i[4], op2_i[2]);
and g260(n415, op2_i[1], op1_i[7]);
and g261(n400, op2_i[4], op1_i[4]);
and g262(n364, op2_i[3], op1_i[6]);
and g263(n331, op2_i[6], op1_i[0], xenc100);
and g264(n386, op2_i[4], op1_i[3]);
and g265(n467, op1_i[5], op2_i[2]);
and g266(n443, op2_i[3], op1_i[4]);
and g267(n406, op2_i[3], op1_i[5]);
and g268(n267, op2_i[4], op1_i[6]);
nand g269(n245, op2_i[5], op1_i[7]);
nand g270(n210, op2_i[7], op1_i[1]);
and g271(n332, op2_i[6], op1_i[1]);
and g272(n343, op2_i[5], op1_i[3]);
and g273(n299, op2_i[3], op1_i[7]);
and g274(n321, op2_i[6], op1_i[3]);
and g275(n273, op2_i[5], op1_i[6]);
and g276(n328, op2_i[6], op1_i[2]);
and g277(n206, op2_i[7], op1_i[2]);
and g278(n357, op2_i[5], op1_i[4]);
and g279(n293, op2_i[6], op1_i[4]);
and g280(n286, op2_i[7], op1_i[3]);
and g281(n262, op2_i[6], op1_i[5]);
and g282(n248, op2_i[6], op1_i[6]);
xnor g283(product_o[6], xenc42, xenc100);
nand g284(n213, op2_i[6], op1_i[0]);
xnor g285(product_o[7], xenc95, xenc117);
nand g286(n211, op2_i[7], op1_i[0]);
and g287(n370, op2_i[4], op1_i[5]);
and g288(n310, op2_i[5], op1_i[5]);
xnor g289(xenc61, n215, n216);
nand g290(n215, op2_i[5], op1_i[0]);
nand g291(n231, op2_i[6], op1_i[7]);
xnor g292(product_o[4], n487, xenc122);
nand g293(n487, op2_i[4], op1_i[0]);
and g294(n279, op2_i[7], op1_i[4]);
and g295(n254, op2_i[7], op1_i[5]);
and g296(n234, op2_i[7], op1_i[6]);
and g297(xenc76, op2_i[0], op1_i[0]);
and g298(xenc98, op2_i[1], op1_i[0]);
and g299(product_o[2], op2_i[2], op1_i[0]);
and g300(product_o[3], op2_i[3], op1_i[0]);
xnor g301(xenc0, n205, keyinput0);
xor g302(xenc1, n281, keyinput1);
xnor g303(xenc2, n268, keyinput2);
xnor g304(xenc3, n469, keyinput3);
xnor g305(xenc4, n315, keyinput4);
xor g306(xenc5, n226, keyinput5);
xnor g307(xenc6, n225, keyinput6);
xnor g308(xenc7, n327, keyinput7);
xor g309(xenc8, n224, keyinput8);
xor g310(xenc9, n317, keyinput9);
xor g311(xenc10, n417, keyinput10);
xor g312(xenc11, n372, keyinput11);
xnor g313(xenc12, n238, keyinput12);
xor g314(xenc13, n433, keyinput13);
xnor g315(xenc14, n297, keyinput14);
xor g316(xenc15, n345, keyinput15);
xor g317(xenc16, n359, keyinput16);
xor g318(xenc17, n435, keyinput17);
xor g319(xenc18, n239, keyinput18);
xnor g320(xenc19, n311, keyinput19);
xnor g321(xenc20, n247, keyinput20);
xnor g322(xenc21, n237, keyinput21);
xnor g323(xenc22, n391, keyinput22);
xor g324(xenc23, n360, keyinput23);
xor g325(xenc24, n404, keyinput24);
xnor g326(xenc25, n368, keyinput25);
xnor g327(xenc26, n248, keyinput26);
xnor g328(xenc27, n446, keyinput27);
xor g329(xenc28, n383, keyinput28);
xor g330(xenc29, n449, keyinput29);
xnor g331(product_o[11], xenc30, keyinput30);
xor g332(xenc31, n409, keyinput31);
xnor g333(xenc32, n382, keyinput32);
xnor g334(xenc33, n380, keyinput33);
xor g335(xenc34, n301, keyinput34);
xor g336(xenc35, n219, keyinput35);
xor g337(xenc36, n437, keyinput36);
xor g338(xenc37, n329, keyinput37);
xor g339(xenc38, n381, keyinput38);
xnor g340(xenc39, n486, keyinput39);
xnor g341(xenc40, n309, keyinput40);
xnor g342(xenc41, n337, keyinput41);
xor g343(xenc42, n213, keyinput42);
xnor g344(xenc43, n374, keyinput43);
xor g345(xenc44, n306, keyinput44);
xnor g346(xenc45, n324, keyinput45);
xor g347(xenc46, n466, keyinput46);
xnor g348(xenc47, n434, keyinput47);
xor g349(xenc48, n259, keyinput48);
xnor g350(xenc49, n477, keyinput49);
xor g351(xenc50, n269, keyinput50);
xor g352(xenc51, n384, keyinput51);
xor g353(xenc52, n304, keyinput52);
xor g354(xenc53, n280, keyinput53);
xor g355(xenc54, n475, keyinput54);
xnor g356(xenc55, n289, keyinput55);
xor g357(xenc56, n314, keyinput56);
xor g358(xenc57, n270, keyinput57);
xnor g359(xenc58, n254, keyinput58);
xnor g360(xenc59, n427, keyinput59);
xor g361(xenc60, n332, keyinput60);
xnor g362(product_o[5], xenc61, keyinput61);
xor g363(xenc62, n233, keyinput62);
xor g364(xenc63, n463, keyinput63);
xor g365(xenc64, n257, keyinput64);
xnor g366(xenc65, n299, keyinput65);
xnor g367(xenc66, n416, keyinput66);
xnor g368(xenc67, n260, keyinput67);
xor g369(xenc68, n326, keyinput68);
xor g370(xenc69, n249, keyinput69);
xor g371(xenc70, n441, keyinput70);
xor g372(xenc71, n261, keyinput71);
xor g373(xenc72, n208, keyinput72);
xnor g374(xenc73, n353, keyinput73);
xor g375(xenc74, n483, keyinput74);
xor g376(xenc75, n385, keyinput75);
xnor g377(product_o[0], xenc76, keyinput76);
xnor g378(xenc77, n232, keyinput77);
xor g379(xenc78, n465, keyinput78);
xor g380(xenc79, n440, keyinput79);
xor g381(xenc80, n295, keyinput80);
xnor g382(xenc81, n476, keyinput81);
xor g383(xenc82, n210, keyinput82);
xnor g384(xenc83, n220, keyinput83);
xnor g385(xenc84, n349, keyinput84);
xnor g386(xenc85, n431, keyinput85);
xnor g387(xenc86, n370, keyinput86);
xor g388(xenc87, n419, keyinput87);
xor g389(product_o[12], xenc88, keyinput88);
xnor g390(xenc89, n398, keyinput89);
xnor g391(xenc90, n338, keyinput90);
xnor g392(xenc91, n438, keyinput91);
xor g393(xenc92, n399, keyinput92);
xor g394(xenc93, n243, keyinput93);
xnor g395(xenc94, n292, keyinput94);
xnor g396(xenc95, n211, keyinput95);
xnor g397(xenc96, n262, keyinput96);
xnor g398(xenc97, n234, keyinput97);
xnor g399(product_o[1], xenc98, keyinput98);
xor g400(xenc99, n401, keyinput99);
xnor g401(xenc100, n214, keyinput100);
xor g402(xenc101, n207, keyinput101);
xor g403(xenc102, n339, keyinput102);
xor g404(xenc103, n462, keyinput103);
xnor g405(xenc104, n396, keyinput104);
xnor g406(xenc105, n356, keyinput105);
xnor g407(xenc106, n267, keyinput106);
xnor g408(xenc107, n390, keyinput107);
xor g409(xenc108, n415, keyinput108);
xnor g410(xenc109, n282, keyinput109);
xnor g411(xenc110, n478, keyinput110);
xnor g412(xenc111, n206, keyinput111);
xnor g413(xenc112, n241, keyinput112);
xor g414(xenc113, n286, keyinput113);
xnor g415(xenc114, n414, keyinput114);
xnor g416(xenc115, n221, keyinput115);
xor g417(xenc116, n316, keyinput116);
xnor g418(xenc117, n212, keyinput117);
xnor g419(xenc118, n358, keyinput118);
xnor g420(xenc119, n387, keyinput119);
xnor g421(xenc120, n285, keyinput120);
xnor g422(xenc121, n278, keyinput121);
xor g423(xenc122, n218, keyinput122);
xor g424(xenc123, n369, keyinput123);
xor g425(xenc124, n305, keyinput124);
xor g426(xenc125, n283, keyinput125);
xor g427(xenc126, n240, keyinput126);
xor g428(xenc127, n418, keyinput127);
endmodule
