library verilog;
use verilog.vl_types.all;
entity xnor_based_carry_lookahead_adder32_tb is
end xnor_based_carry_lookahead_adder32_tb;
