// Verilog File 
module equal_segmentation_adder32_ant_enc32.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput1,keyinput0,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,result_o[0],
result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],result_o[7],result_o[8],result_o[9],result_o[10],
result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],result_o[17],result_o[18],result_o[19],result_o[20],
result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],result_o[27],result_o[28],result_o[29],result_o[30],
result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput1,keyinput0,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n76, n77, n78, n81, n82, n85, n86, n89, n90, 
n93, n94, n101, n102, n105, n106, n97, n98, n109, n110, 
n116, n117, n120, n121, n124, n125, n128, n130, n131, n134, 
n135, n138, n139, n142, n143, n113, n146, n147, n151, n152, 
n155, n157, n158, n161, n162, n165, n166, n169, n170, n173, 
n174, n177, n178, n129, n148, n181, n156, n79, n80, n159, 
n160, n132, n133, n122, n123, n95, n96, n175, n176, n149, 
n150, n118, n119, n91, n92, n171, n172, n144, n145, n103_ant0, 
n104, n103, n114, n115, n87, n88, n167, n168, n140, n141, 
n107, n108, n83, n84, n163, n164, n136, n137, n126, n127, 
n111, n112, n179, n180, n153, n154, n99, n100, antisat_out, in0xor_0, 
in1xor_0, inter30_0, in2xor_0, in3xor_0, inter29_0, in4xor_0, in5xor_0, inter28_0, in6xor_0, in7xor_0, 
inter27_0, in8xor_0, in9xor_0, inter26_0, in10xor_0, in11xor_0, inter25_0, in12xor_0, in13xor_0, inter24_0, 
in14xor_0, in15xor_0, inter23_0, in16xor_0, in17xor_0, inter22_0, in18xor_0, in19xor_0, inter21_0, in20xor_0, 
in21xor_0, inter20_0, in22xor_0, in23xor_0, inter19_0, in24xor_0, in25xor_0, inter18_0, in26xor_0, in27xor_0, 
inter17_0, in28xor_0, in29xor_0, inter16_0, in30xor_0, in31xor_0, inter15_0, inter14_0, inter13_0, inter12_0, 
inter11_0, inter10_0, inter9_0, inter8_0, inter7_0, inter6_0, inter5_0, inter4_0, inter3_0, inter2_0, 
inter1_0, antisat_g_0, in0xor_b_0, in1xor_b_0, inter30_b_0, in2xor_b_0, in3xor_b_0, inter29_b_0, in4xor_b_0, in5xor_b_0, 
inter28_b_0, in6xor_b_0, in7xor_b_0, inter27_b_0, in8xor_b_0, in9xor_b_0, inter26_b_0, in10xor_b_0, in11xor_b_0, inter25_b_0, 
in12xor_b_0, in13xor_b_0, inter24_b_0, in14xor_b_0, in15xor_b_0, inter23_b_0, in16xor_b_0, in17xor_b_0, inter22_b_0, in18xor_b_0, 
in19xor_b_0, inter21_b_0, in20xor_b_0, in21xor_b_0, inter20_b_0, in22xor_b_0, in23xor_b_0, inter19_b_0, in24xor_b_0, in25xor_b_0, 
inter18_b_0, in26xor_b_0, in27xor_b_0, inter17_b_0, in28xor_b_0, in29xor_b_0, inter16_b_0, in30xor_b_0, in31xor_b_0, inter15_b_0, 
inter14_b_0, inter13_b_0, inter12_b_0, inter11_b_0, inter10_b_0, inter9_b_0, inter8_b_0, inter7_b_0, inter6_b_0, inter5_b_0, 
inter4_b_0, inter3_b_0, inter2_b_0, inter1_b_0, inter0_b_0, antisat_gbar_0;

xor g0(result_o[9], add2_i[9], n76);
xor g1(result_o[8], add2_i[8], add1_i[8]);
xor g2(result_o[7], n77, n78);
xor g3(n78, add2_i[7], add1_i[7]);
xor g4(result_o[6], add2_i[6], n81);
xor g5(n81, n82, add1_i[6]);
xor g6(result_o[5], add2_i[5], n85);
xor g7(n85, n86, add1_i[5]);
xor g8(result_o[4], add2_i[4], n89);
xor g9(n89, n90, add1_i[4]);
xor g10(result_o[3], add2_i[3], n93);
xor g11(n93, n94, add1_i[3]);
xor g12(result_o[31], add2_i[31], n101);
xor g13(n101, n102, add1_i[31]);
xor g14(result_o[30], add2_i[30], n105);
xor g15(n105, n106, add1_i[30]);
xor g16(result_o[2], add2_i[2], n97);
xor g17(n97, n98, add1_i[2]);
xor g18(result_o[29], add2_i[29], n109);
xor g19(n109, n110, add1_i[29]);
xor g20(result_o[28], add2_i[28], n116);
xor g21(n116, n117, add1_i[28]);
xor g22(result_o[27], add2_i[27], n120);
xor g23(n120, n121, add1_i[27]);
xor g24(result_o[26], add2_i[26], n124);
xor g25(n124, n125, add1_i[26]);
xor g26(result_o[25], add2_i[25], n128);
xor g27(result_o[24], add2_i[24], add1_i[24]);
xor g28(result_o[23], n130, n131);
xor g29(n131, add2_i[23], add1_i[23]);
xor g30(result_o[22], add2_i[22], n134);
xor g31(n134, n135, add1_i[22]);
xor g32(result_o[21], add2_i[21], n138);
xor g33(n138, n139, add1_i[21]);
xor g34(result_o[20], add2_i[20], n142);
xor g35(n142, n143, add1_i[20]);
xor g36(result_o[1], add2_i[1], n113);
xor g37(result_o[19], add2_i[19], n146);
xor g38(n146, n147, add1_i[19]);
xor g39(result_o[18], add2_i[18], n151);
xor g40(n151, n152, add1_i[18]);
xor g41(result_o[17], add2_i[17], n155);
xor g42(result_o[16], add2_i[16], add1_i[16]);
xor g43(result_o[15], n157, n158);
xor g44(n158, add2_i[15], add1_i[15]);
xor g45(result_o[14], add2_i[14], n161);
xor g46(n161, n162, add1_i[14]);
xor g47(result_o[13], add2_i[13], n165);
xor g48(n165, n166, add1_i[13]);
xor g49(result_o[12], add2_i[12], n169);
xor g50(n169, n170, add1_i[12]);
xor g51(result_o[11], add2_i[11], n173);
xor g52(n173, n174, add1_i[11]);
xor g53(result_o[10], add2_i[10], n177);
xor g54(n177, n178, add1_i[10]);
xor g55(result_o[0], add2_i[0], add1_i[0]);
xnor g56(n128, n129, add1_i[25]);
nand g57(n129, add2_i[24], add1_i[24]);
xnor g58(n113, n148, add1_i[1]);
nand g59(n148, add2_i[0], add1_i[0]);
xnor g60(n76, n181, add1_i[9]);
nand g61(n181, add2_i[8], add1_i[8]);
xnor g62(n155, n156, add1_i[17]);
nand g63(n156, add2_i[16], add1_i[16]);
nand g64(n77, n79, n80);
nand g65(n79, add1_i[6], n82);
nand g66(n157, n159, n160);
nand g67(n159, add1_i[14], n162);
nand g68(n130, n132, n133);
nand g69(n132, add1_i[22], n135);
nand g70(n121, n122, n123);
nand g71(n122, add1_i[26], n125);
nand g72(n123, add2_i[26], n124);
nand g73(n94, n95, n96);
nand g74(n95, add1_i[2], n98);
nand g75(n96, add2_i[2], n97);
nand g76(n174, n175, n176);
nand g77(n175, add1_i[10], n178);
nand g78(n176, add2_i[10], n177);
nand g79(n147, n149, n150);
nand g80(n149, add1_i[18], n152);
nand g81(n150, add2_i[18], n151);
nand g82(n117, n118, n119);
nand g83(n118, add1_i[27], n121);
nand g84(n119, add2_i[27], n120);
nand g85(n90, n91, n92);
nand g86(n91, add1_i[3], n94);
nand g87(n92, add2_i[3], n93);
nand g88(n170, n171, n172);
nand g89(n171, add1_i[11], n174);
nand g90(n172, add2_i[11], n173);
nand g91(n143, n144, n145);
nand g92(n144, add1_i[19], n147);
nand g93(n145, add2_i[19], n146);
nand g94(n102, n103_ant0, n104);
nand g95(n103, add1_i[30], n106);
nand g96(n104, add2_i[30], n105);
nand g97(n110, n114, n115);
nand g98(n114, add1_i[28], n117);
nand g99(n115, add2_i[28], n116);
nand g100(n86, n87, n88);
nand g101(n87, add1_i[4], n90);
nand g102(n88, add2_i[4], n89);
nand g103(n166, n167, n168);
nand g104(n167, add1_i[12], n170);
nand g105(n168, add2_i[12], n169);
nand g106(n139, n140, n141);
nand g107(n140, add1_i[20], n143);
nand g108(n141, add2_i[20], n142);
nand g109(n106, n107, n108);
nand g110(n107, add1_i[29], n110);
nand g111(n108, add2_i[29], n109);
nand g112(n82, n83, n84);
nand g113(n83, add1_i[5], n86);
nand g114(n84, add2_i[5], n85);
nand g115(n162, n163, n164);
nand g116(n163, add1_i[13], n166);
nand g117(n164, add2_i[13], n165);
nand g118(n135, n136, n137);
nand g119(n136, add1_i[21], n139);
nand g120(n137, add2_i[21], n138);
nand g121(n80, add2_i[6], n81);
nand g122(n160, add2_i[14], n161);
nand g123(n133, add2_i[22], n134);
nand g124(n125, n126, n127);
nand g125(n127, add1_i[25], add1_i[24], add2_i[24]);
nand g126(n126, add2_i[25], n128);
nand g127(n98, n111, n112);
nand g128(n112, add1_i[1], add1_i[0], add2_i[0]);
nand g129(n111, add2_i[1], n113);
nand g130(n178, n179, n180);
nand g131(n180, add2_i[8], add1_i[8], add1_i[9]);
nand g132(n179, add2_i[9], n76);
nand g133(n152, n153, n154);
nand g134(n154, add1_i[17], add1_i[16], add2_i[16]);
nand g135(n153, add2_i[17], n155);
nand g136(result_o[32], n99, n100);
nand g137(n99, add1_i[31], n102);
nand g138(n100, add2_i[31], n101);
xor g139(n103_ant0, n103, antisat_out);
and g140(inter30_0, in0xor_0, in1xor_0);
and g141(inter29_0, in2xor_0, in3xor_0);
and g142(inter28_0, in4xor_0, in5xor_0);
and g143(inter27_0, in6xor_0, in7xor_0);
and g144(inter26_0, in8xor_0, in9xor_0);
and g145(inter25_0, in10xor_0, in11xor_0);
and g146(inter24_0, in12xor_0, in13xor_0);
and g147(inter23_0, in14xor_0, in15xor_0);
and g148(inter22_0, in16xor_0, in17xor_0);
and g149(inter21_0, in18xor_0, in19xor_0);
and g150(inter20_0, in20xor_0, in21xor_0);
and g151(inter19_0, in22xor_0, in23xor_0);
and g152(inter18_0, in24xor_0, in25xor_0);
and g153(inter17_0, in26xor_0, in27xor_0);
and g154(inter16_0, in28xor_0, in29xor_0);
and g155(inter15_0, in30xor_0, in31xor_0);
and g156(inter14_0, inter30_0, inter29_0);
and g157(inter13_0, inter28_0, inter27_0);
and g158(inter12_0, inter26_0, inter25_0);
and g159(inter11_0, inter24_0, inter23_0);
and g160(inter10_0, inter22_0, inter21_0);
and g161(inter9_0, inter20_0, inter19_0);
and g162(inter8_0, inter18_0, inter17_0);
and g163(inter7_0, inter16_0, inter15_0);
and g164(inter6_0, inter14_0, inter13_0);
and g165(inter5_0, inter12_0, inter11_0);
and g166(inter4_0, inter10_0, inter9_0);
and g167(inter3_0, inter8_0, inter7_0);
and g168(inter2_0, inter6_0, inter5_0);
and g169(inter1_0, inter4_0, inter3_0);
and g170(antisat_g_0, inter2_0, inter1_0);
xor g171(in0xor_0, n128, keyinput0);
xor g172(in1xor_0, n121, keyinput1);
xor g173(in2xor_0, n107, keyinput2);
xor g174(in3xor_0, n108, keyinput3);
xor g175(in4xor_0, n123, keyinput4);
xor g176(in5xor_0, n124, keyinput5);
xor g177(in6xor_0, n126, keyinput6);
xor g178(in7xor_0, n109, keyinput7);
xor g179(in8xor_0, add2_i[26], keyinput8);
xor g180(in9xor_0, n116, keyinput9);
xor g181(in10xor_0, add1_i[25], keyinput10);
xor g182(in11xor_0, n127, keyinput11);
xor g183(in12xor_0, add2_i[27], keyinput12);
xor g184(in13xor_0, n129, keyinput13);
xor g185(in14xor_0, add2_i[25], keyinput14);
xor g186(in15xor_0, add1_i[26], keyinput15);
xor g187(in16xor_0, n110, keyinput16);
xor g188(in17xor_0, add2_i[28], keyinput17);
xor g189(in18xor_0, add1_i[24], keyinput18);
xor g190(in19xor_0, add2_i[29], keyinput19);
xor g191(in20xor_0, n119, keyinput20);
xor g192(in21xor_0, add1_i[28], keyinput21);
xor g193(in22xor_0, n120, keyinput22);
xor g194(in23xor_0, add1_i[29], keyinput23);
xor g195(in24xor_0, add2_i[24], keyinput24);
xor g196(in25xor_0, add1_i[30], keyinput25);
xor g197(in26xor_0, n118, keyinput26);
xor g198(in27xor_0, add1_i[27], keyinput27);
xor g199(in28xor_0, n117, keyinput28);
xor g200(in29xor_0, n106, keyinput29);
xor g201(in30xor_0, n114, keyinput30);
xor g202(in31xor_0, n115, keyinput31);
and g203(inter30_b_0, in0xor_b_0, in1xor_b_0);
and g204(inter29_b_0, in2xor_b_0, in3xor_b_0);
and g205(inter28_b_0, in4xor_b_0, in5xor_b_0);
and g206(inter27_b_0, in6xor_b_0, in7xor_b_0);
and g207(inter26_b_0, in8xor_b_0, in9xor_b_0);
and g208(inter25_b_0, in10xor_b_0, in11xor_b_0);
and g209(inter24_b_0, in12xor_b_0, in13xor_b_0);
and g210(inter23_b_0, in14xor_b_0, in15xor_b_0);
and g211(inter22_b_0, in16xor_b_0, in17xor_b_0);
and g212(inter21_b_0, in18xor_b_0, in19xor_b_0);
and g213(inter20_b_0, in20xor_b_0, in21xor_b_0);
and g214(inter19_b_0, in22xor_b_0, in23xor_b_0);
and g215(inter18_b_0, in24xor_b_0, in25xor_b_0);
and g216(inter17_b_0, in26xor_b_0, in27xor_b_0);
and g217(inter16_b_0, in28xor_b_0, in29xor_b_0);
and g218(inter15_b_0, in30xor_b_0, in31xor_b_0);
and g219(inter14_b_0, inter30_b_0, inter29_b_0);
and g220(inter13_b_0, inter28_b_0, inter27_b_0);
and g221(inter12_b_0, inter26_b_0, inter25_b_0);
and g222(inter11_b_0, inter24_b_0, inter23_b_0);
and g223(inter10_b_0, inter22_b_0, inter21_b_0);
and g224(inter9_b_0, inter20_b_0, inter19_b_0);
and g225(inter8_b_0, inter18_b_0, inter17_b_0);
and g226(inter7_b_0, inter16_b_0, inter15_b_0);
and g227(inter6_b_0, inter14_b_0, inter13_b_0);
and g228(inter5_b_0, inter12_b_0, inter11_b_0);
and g229(inter4_b_0, inter10_b_0, inter9_b_0);
and g230(inter3_b_0, inter8_b_0, inter7_b_0);
and g231(inter2_b_0, inter6_b_0, inter5_b_0);
and g232(inter1_b_0, inter4_b_0, inter3_b_0);
and g233(inter0_b_0, inter2_b_0, inter1_b_0);
xor g234(in0xor_b_0, n128, keyinput32);
xor g235(in1xor_b_0, n121, keyinput33);
xor g236(in2xor_b_0, n107, keyinput34);
xor g237(in3xor_b_0, n108, keyinput35);
xor g238(in4xor_b_0, n123, keyinput36);
xor g239(in5xor_b_0, n124, keyinput37);
xor g240(in6xor_b_0, n126, keyinput38);
xor g241(in7xor_b_0, n109, keyinput39);
xor g242(in8xor_b_0, add2_i[26], keyinput40);
xor g243(in9xor_b_0, n116, keyinput41);
xor g244(in10xor_b_0, add1_i[25], keyinput42);
xor g245(in11xor_b_0, n127, keyinput43);
xor g246(in12xor_b_0, add2_i[27], keyinput44);
xor g247(in13xor_b_0, n129, keyinput45);
xor g248(in14xor_b_0, add2_i[25], keyinput46);
xor g249(in15xor_b_0, add1_i[26], keyinput47);
xor g250(in16xor_b_0, n110, keyinput48);
xor g251(in17xor_b_0, add2_i[28], keyinput49);
xor g252(in18xor_b_0, add1_i[24], keyinput50);
xor g253(in19xor_b_0, add2_i[29], keyinput51);
xor g254(in20xor_b_0, n119, keyinput52);
xor g255(in21xor_b_0, add1_i[28], keyinput53);
xor g256(in22xor_b_0, n120, keyinput54);
xor g257(in23xor_b_0, add1_i[29], keyinput55);
xor g258(in24xor_b_0, add2_i[24], keyinput56);
xor g259(in25xor_b_0, add1_i[30], keyinput57);
xor g260(in26xor_b_0, n118, keyinput58);
xor g261(in27xor_b_0, add1_i[27], keyinput59);
xor g262(in28xor_b_0, n117, keyinput60);
xor g263(in29xor_b_0, n106, keyinput61);
xor g264(in30xor_b_0, n114, keyinput62);
xor g265(in31xor_b_0, n115, keyinput63);
not g266(antisat_gbar_0, inter0_b_0);
and g267(antisat_out, antisat_g_0, antisat_gbar_0);
endmodule
