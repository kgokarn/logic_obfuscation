// Verilog File 
module underdesigned_multiplier8_aor_enc128.bench (op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,product_o[0],product_o[1],product_o[2],product_o[3],product_o[4],
product_o[5],product_o[6],product_o[7],product_o[8],product_o[9],product_o[10],product_o[11],product_o[12],product_o[13],product_o[14],
product_o[15]);

input op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127;


output product_o[0], product_o[1], product_o[2], product_o[3], product_o[4], product_o[5], product_o[6], product_o[7], product_o[8], 
product_o[9], product_o[10], product_o[11], product_o[12], product_o[13], product_o[14], product_o[15];

wire n158, n159, n160, n161, xenc81, xenc119, n163, n171, n170, 
xenc127, n174, xenc0, xenc61, n186, n187, n183, xenc42, xenc53, n232, 
n229, xenc89, n221, xenc115, n235, n274, xenc86, n272, n298, xenc124, 
n268, n320, n319, n169, n332, n333, n327, xenc24, n334, n335, 
n331, n336, n337, n329, xenc97, n341, n338, xenc122, xenc33, n343, 
xenc110, n351, n352, n353, n347, n354, n355, n356, xenc19, n380, 
n381, n382, n383, n378, xenc9, xenc102, xenc85, n396, n391, n368, 
n392, n389, n415, n416, n385, xenc67, xenc44, n386, n289, n288, 
n312, n303, xenc52, n309, n456, n457, n455, n462, n435, n417, 
xenc3, n441, n420, xenc25, n244, n215, xenc78, n245, n243, n246, 
n278, n276, n277, n280, n279, n478, xenc18, xenc77, xenc99, n479, 
xenc106, n283, n284, n282, n247, xenc107, n316, n374, n149, n167, 
xenc27, xenc39, n195, n143, n480, xenc114, xenc65, n162, n166, n318, 
xenc116, n317, n315, n192, n193, n184, n372, n373, n216, n249, 
n250, xenc38, xenc96, n481, xenc41, xenc29, xenc83, n418, n348, n349, 
n342, n164, xenc51, n286, xenc40, n251, n148, n377, n313, n447, 
n448, n419, xenc48, n449, xenc22, n445, n294, n444, n446, xenc91, 
n292, n275, xenc47, n296, n291, n293, n285, n287, xenc31, n345, 
n344, xenc80, xenc57, n214, n212, n213, xenc82, n376, n150, n375, 
xenc126, n431, n182, n197, n194, xenc100, n199, xenc5, n311, n314, 
xenc79, n200, n228, n145, xenc120, n191, xenc28, n147, n270, n271, 
n222, xenc12, xenc16, n482, xenc74, xenc26, n225, n227, n226, n483, 
xenc66, xenc14, n231, n233, xenc88, n201, n198, n346, xenc1, n442, 
n470, xenc73, xenc36, n422, n153, n409, n155, n402, n151, n157, 
n460, n452, n154, n152, n425, n304, xenc37, xenc34, xenc98, n371, 
n369, n454, n414, xenc50, n384, n297, xenc109, xenc17, n269, n458, 
xenc105, xenc11, n453, n451, xenc84, n406, xenc15, n400, n393, xenc113, 
n379, xenc93, n394, n395, xenc46, n404, n403, n405, xenc4, xenc43, 
n267, n310, xenc32, n305, xenc70, n308, n306, n307, n484, xenc55, 
xenc6, n472, n471, n473, xenc64, xenc59, n397, n399, n398, xenc49, 
n181, xenc117, n180, n263, xenc118, n437, n436, n255, n242, n156, 
n321, n325, n210, n209, n236, n323, n324, n175, xenc56, n241, 
n252, n230, xenc76, n240, n421, n290, n273, n330, xenc30, n328, 
n172, xenc108, n177, n322, n430, xenc35, n211, n220, n144, n339, 
n190, n189, n461, xenc94, n439, n438, xenc123, n440, n432, xenc111, 
n295, n434, n433, n358, n359, n360, n258, n259, xenc104, n260, 
n361, xenc103, n363, n362, n387, xenc112, xenc92, n388, n390, xenc45, 
xenc69, n234, n264, n266, n265, n218, xenc121, n219, n188, n204, 
n205, xenc58, xenc2, n206, n463, n464, xenc60, n465, n299, n300, 
n261, n301, n237, n238, n208, n239, n207, n173, xenc20, xenc13, 
n411, n401, n410, n407, n408, n146, xenc71, xenc87, n350, n485, 
n443, n370, xenc75, xenc23, n366, n367, xenc21, n469, n450, n468, 
xenc95, xenc62, n256, n257, n262, n476, n477, n466, n467, xenc54, 
n365, n326, n364, xenc10, n429, n428, xenc7, xenc90, n302, n423, 
n424, n253, xenc72, n254, n426, xenc68, n427, n340, n412, n413, 
n357, n223, n224, xenc8, n475, n474, n202, xenc125, n203, n486, 
xenc63, n178, xenc101, n179;

xor g0(product_o[9], n158, n159);
xor g1(xenc81, n160, n161);
xor g2(n160, xenc119, n163);
xor g3(xenc127, n171, n170);
xor g4(xenc61, n174, xenc0);
xor g5(n183, n186, n187);
xor g6(n232, xenc42, xenc53);
xor g7(n221, n229, xenc89);
xor g8(n229, xenc115, n235);
xor g9(n272, n274, xenc86);
xor g10(n268, n298, xenc124);
xor g11(n169, n320, n319);
xor g12(n320, n332, n333);
xor g13(n170, n327, xenc24);
xor g14(n331, n334, n335);
xor g15(n329, n336, n337);
xor g16(n338, xenc97, n341);
xor g17(n343, xenc122, xenc33);
xor g18(n332, xenc110, n351);
xor g19(n347, n352, n353);
xor g20(n335, n354, n355);
xor g21(n354, n356, xenc19);
xor g22(n352, n380, n381);
xor g23(n381, n382, n383);
xor g24(n353, n378, xenc9);
xor g25(n159, xenc102, xenc85);
xor g26(n368, n396, n391);
xor g27(n396, n392, n389);
xor g28(n385, n415, n416);
xor g29(n386, xenc67, xenc44);
xor g30(n312, n289, n288);
xor g31(n309, n303, xenc52);
xor g32(n455, n456, n457);
xor g33(n417, n462, n435);
xor g34(n420, xenc3, n441);
nand g35(n215, xenc25, n244);
nand g36(n243, xenc78, n245);
nand g37(n244, n245, n246);
and g38(n278, n159, n158);
nand g39(n246, n276, n277);
nand g40(n276, n280, n279);
nand g41(n277, n278, n279);
xnor g42(xenc18, n478, n279);
nor g43(n478, n278, n280);
xnor g44(xenc99, xenc77, n245);
nor g45(n479, n246, xenc78);
nor g46(n279, xenc78, xenc106);
and g47(n282, n283, n284);
nor g48(n247, n284, n283);
nand g49(n316, n353, n352, xenc107);
not g50(n149, n374);
nand g51(n167, n319, n320);
xnor g52(product_o[13], xenc27, xenc39);
nor g53(n480, n195, n143);
nand g54(n162, xenc114, xenc65);
nand g55(n318, n166, n167);
nand g56(n158, xenc116, n316);
nand g57(n315, n163, n317);
nand g58(n317, n161, xenc119);
nand g59(n184, n192, n193);
nand g60(n192, n143, xenc39);
nand g61(n193, xenc39, n195);
and g62(n163, n316, n372);
nand g63(n372, n373, n374);
nand g64(n373, n353, n352);
nor g65(n245, n216, n249);
and g66(n249, n250, xenc38);
nor g67(n216, xenc38, n250);
xnor g68(n250, xenc96, n221);
nor g69(n280, xenc85, xenc102);
xor g70(xenc41, xenc114, n481);
nand g71(n481, n166, n167);
xnor g72(n418, xenc29, xenc83);
xnor g73(n333, n348, n349);
nand g74(n348, n335, n334);
xnor g75(n164, n342, n343);
nand g76(n342, n332, n333);
xnor g77(n286, n272, xenc51);
nand g78(n166, n170, n169, n171);
nand g79(n251, n289, n288, xenc40);
not g80(n148, n286);
nand g81(n313, xenc9, n378, n377);
nand g82(n419, n447, n448);
or g83(n447, n382, n383);
nand g84(n448, n380, xenc48);
nand g85(n449, n383, n382);
nand g86(n294, xenc22, n445);
or g87(n444, xenc83, xenc67);
nand g88(n445, n446, xenc29);
nand g89(n446, xenc67, xenc83);
nand g90(n275, xenc91, n292);
nand g91(n291, xenc47, n296);
nand g92(n292, n293, n294);
or g93(n293, xenc47, n296);
nand g94(n283, xenc38, n285);
nand g95(n285, n286, n287);
nand g96(n287, n288, n289);
and g97(n161, xenc31, n345);
nand g98(n344, xenc122, xenc33);
nand g99(n345, n332, n333, n343);
nand g100(n195, xenc80, xenc57);
nand g101(n212, n216, n214);
nand g102(n213, n214, n215);
nand g103(n374, xenc85, xenc82);
nand g104(n375, n376, n150);
nand g105(n376, n378, xenc9);
not g106(n150, n377);
xnor g107(n289, xenc126, xenc47);
xnor g108(n431, n294, n296);
nor g109(n194, n182, n197);
and g110(n197, xenc100, n199);
nor g111(n182, n199, xenc100);
xnor g112(n314, xenc5, n311);
nand g113(n200, n229, xenc89, xenc79);
not g114(n145, n228);
nand g115(n191, n235, xenc115, xenc120);
not g116(n147, xenc28);
nand g117(n222, n270, n271);
nand g118(n270, n274, xenc86);
nand g119(n271, n272, xenc51);
xnor g120(xenc16, xenc12, n169);
nand g121(n482, n170, n171);
nand g122(n225, xenc74, xenc26);
nand g123(n226, n227, n228);
nand g124(n227, n229, xenc89);
nand g125(n284, n311, xenc5);
xnor g126(product_o[12], n483, n214);
nor g127(n483, n215, n216);
nand g128(n228, n191, xenc66);
nand g129(n231, xenc28, xenc14);
nand g130(n233, xenc115, n235);
not g131(n143, xenc88);
and g132(n319, n327, xenc24);
and g133(n198, xenc74, n201);
and g134(n346, n349, n334, n335);
xnor g135(n470, xenc1, n442);
xnor g136(n422, xenc73, xenc36);
nor g137(n402, n153, n409, n155);
nor g138(n452, n151, n157, n460);
nor g139(n304, n154, n152, n425);
nor g140(n311, n386, n385);
xnor g141(n349, xenc37, xenc34);
xnor g142(n369, xenc98, n371);
xnor g143(n383, n454, n455);
xnor g144(n337, n409, n414);
nor g145(n414, n153, n155);
nor g146(n377, n311, xenc50);
and g147(n384, n385, n386);
xnor g148(n274, n297, xenc109);
xnor g149(n297, xenc17, n269);
nor g150(n458, n155, n152);
xnor g151(n380, xenc105, xenc11);
xnor g152(n451, n452, n453);
xnor g153(n355, xenc84, n406);
xnor g154(n406, xenc15, n400);
nand g155(n379, n393, xenc113);
or g156(n393, xenc98, n371);
nand g157(n394, xenc37, xenc93);
nand g158(n395, n371, xenc98);
and g159(n371, xenc46, n404);
or g160(n403, n356, xenc19);
nand g161(n404, n355, n405);
nand g162(n405, xenc19, n356);
nand g163(n267, xenc4, xenc43);
or g164(n305, n310, xenc32);
nand g165(n306, xenc70, n308);
nand g166(n307, xenc32, n310);
xnor g167(product_o[14], n484, xenc55);
nor g168(n484, n184, n182);
nand g169(n441, xenc6, n472);
or g170(n471, n456, n454);
nand g171(n472, n473, n457);
nand g172(n473, n454, n456);
and g173(n391, xenc64, xenc59);
nand g174(n397, xenc15, xenc84);
nand g175(n398, n399, n400);
or g176(n399, xenc84, xenc15);
nand g177(xenc117, xenc49, n181);
nand g178(n181, n182, xenc55);
nand g179(n180, xenc55, n184);
xnor g180(n298, n263, xenc118);
xnor g181(n462, n437, n436);
nor g182(n242, n151, n155, n255);
nor g183(n325, n153, n156, n321);
xnor g184(n236, n210, n209);
xnor g185(n175, n323, n324);
xnor g186(n324, n325, xenc56);
xnor g187(n230, n241, n252);
xnor g188(n252, xenc76, n240);
xnor g189(n288, n421, xenc32);
xnor g190(n421, n310, n308);
xnor g191(n273, n255, n290);
nor g192(n290, n155, n151);
nor g193(n327, n330, xenc30);
nor g194(n172, n327, n328);
and g195(n328, xenc30, n330);
xnor g196(n177, n321, xenc108);
nor g197(n322, n156, n153);
xnor g198(n416, n425, n430);
nor g199(n430, n152, n154);
nand g200(n211, n221, xenc96, xenc35);
not g201(n144, n220);
xnor g202(n330, n338, n339);
xnor g203(n199, n190, n189);
xnor g204(n351, n460, n461);
nor g205(n461, n157, n151);
nand g206(n296, xenc94, n439);
or g207(n438, xenc1, n442);
nand g208(n439, xenc123, n441);
nand g209(n440, n442, xenc1);
nand g210(n295, n432, xenc111);
or g211(n432, n437, n436);
nand g212(n433, n434, n435);
nand g213(n434, n436, n437);
nand g214(n334, n358, n359);
or g215(n358, xenc97, n339);
nand g216(n359, n341, n360);
nand g217(n360, n339, xenc97);
nand g218(n235, n258, n259);
or g219(n258, xenc118, n263);
nand g220(n259, xenc104, xenc124);
nand g221(n260, xenc118, n263);
and g222(n339, n361, xenc103);
nand g223(n361, n325, n323);
nand g224(n362, n363, xenc56);
or g225(n363, n323, n325);
nand g226(n378, n387, xenc112);
or g227(n387, n392, n391);
nand g228(n388, n389, xenc92);
nand g229(n390, n391, n392);
nand g230(n234, xenc45, xenc69);
or g231(n264, n269, xenc109);
nand g232(n265, n266, xenc17);
nand g233(n266, xenc109, n269);
and g234(n214, xenc88, n218);
nand g235(n218, xenc121, n220);
nand g236(n219, n221, xenc96);
nor g237(n188, n189, n190);
nand g238(n190, n204, n191);
nand g239(n204, n205, xenc58);
or g240(n205, n210, n209);
nand g241(n206, xenc2, xenc53);
nand g242(n382, n351, xenc110);
nand g243(n435, n463, n464);
nand g244(n463, n452, xenc105);
nand g245(n464, xenc60, n453);
or g246(n465, xenc105, n452);
nand g247(n261, n299, n300);
nand g248(n299, xenc73, n303);
nand g249(n300, n301, xenc36);
or g250(n301, n303, xenc73);
nand g251(n208, n237, n238);
nand g252(n237, xenc76, n241);
nand g253(n238, n239, n240);
or g254(n239, n241, xenc76);
and g255(n171, n172, xenc0, n174);
or g256(n201, n151, n154, n225);
nand g257(n207, n209, n210);
xnor g258(product_o[4], n172, n173);
nand g259(n173, n174, xenc0);
nor g260(product_o[0], n153, n157);
not g261(n153, op1_i[0]);
not g262(n155, op2_i[4]);
nand g263(n356, op1_i[4], n337, op2_i[0]);
nand g264(n456, op1_i[4], op2_i[2], xenc20);
nand g265(n401, xenc13, n411);
nand g266(n410, op2_i[4], op1_i[1]);
nand g267(n411, op1_i[0], op2_i[5]);
not g268(n152, op1_i[2]);
nand g269(n400, n407, n408);
nand g270(n407, op2_i[2], op1_i[3]);
nand g271(n408, op1_i[2], op2_i[3]);
nand g272(n409, op2_i[2], op1_i[2]);
nand g273(n460, op2_i[6], op1_i[0]);
nand g274(n425, op1_i[4], op2_i[4]);
nand g275(n186, op1_i[7], op2_i[7]);
nor g276(n187, n146, xenc71);
not g277(n146, n191);
xnor g278(n350, xenc20, xenc87);
nand g279(n485, op2_i[2], op1_i[4]);
nand g280(n415, op1_i[6], op2_i[2]);
nand g281(n336, op2_i[0], op1_i[4]);
not g282(n151, op1_i[6]);
nand g283(n310, op2_i[2], n416, op1_i[6]);
nand g284(n269, op1_i[7], op2_i[3]);
nand g285(n443, op2_i[5], op1_i[3]);
nand g286(n437, op2_i[7], op1_i[1]);
nand g287(n370, op2_i[1], op1_i[5]);
nand g288(n210, op2_i[7], op1_i[5]);
nand g289(n323, xenc75, xenc23);
nand g290(n366, op2_i[2], op1_i[1]);
nand g291(n367, op1_i[0], op2_i[3]);
nand g292(n450, xenc21, n469);
nand g293(n468, op2_i[6], op1_i[1]);
nand g294(n469, op2_i[7], op1_i[0]);
nand g295(n241, xenc95, xenc62);
nand g296(n256, op2_i[6], op1_i[5]);
nand g297(n257, op2_i[7], op1_i[4]);
nand g298(n262, op2_i[7], op1_i[3]);
nand g299(n263, op1_i[5], op2_i[5]);
nand g300(n442, op1_i[5], op2_i[3]);
nand g301(n436, op1_i[7], op2_i[1]);
nand g302(n209, op1_i[7], op2_i[5]);
not g303(n154, op2_i[6]);
not g304(n157, op2_i[0]);
and g305(n454, n476, n477);
nand g306(n476, op2_i[4], op1_i[3]);
nand g307(n477, op1_i[2], op2_i[5]);
nand g308(n453, n466, n467);
nand g309(n466, op1_i[7], op2_i[0]);
nand g310(n467, op1_i[6], op2_i[1]);
nand g311(n326, xenc54, n365);
nand g312(n364, op2_i[0], op1_i[3]);
nand g313(n365, op2_i[1], op1_i[2]);
nand g314(n308, xenc10, n429);
nand g315(n428, op1_i[7], op2_i[2]);
nand g316(n429, op1_i[6], op2_i[3]);
nand g317(n302, xenc7, xenc90);
nand g318(n423, op2_i[6], op1_i[3]);
nand g319(n424, op2_i[7], op1_i[2]);
nand g320(n240, n253, xenc72);
nand g321(n253, op1_i[7], op2_i[4]);
nand g322(n254, op1_i[6], op2_i[5]);
nand g323(n303, n426, xenc68);
nand g324(n426, op1_i[5], op2_i[4]);
nand g325(n427, op1_i[4], op2_i[5]);
nand g326(n340, op1_i[1], op2_i[3]);
nand g327(n392, op2_i[5], op1_i[1]);
nand g328(n321, op2_i[0], op1_i[2]);
nand g329(n255, op2_i[6], op1_i[4]);
and g330(n357, n412, n413);
nand g331(n412, op2_i[0], op1_i[5]);
nand g332(n413, op1_i[4], op2_i[1]);
nand g333(n220, n201, n223);
nand g334(n223, n224, n225);
nand g335(n224, op1_i[6], op2_i[6]);
and g336(n174, op1_i[1], n177, op2_i[1]);
and g337(n389, op2_i[3], op1_i[3]);
and g338(n341, op2_i[1], op1_i[3]);
not g339(n156, op2_i[2]);
nand g340(n457, xenc8, n475);
nand g341(n474, op1_i[5], op2_i[2]);
nand g342(n475, op1_i[4], op2_i[3]);
and g343(n189, n202, xenc125);
nand g344(n202, op1_i[7], op2_i[6]);
nand g345(n203, op2_i[7], op1_i[6]);
xnor g346(xenc63, n486, n177);
nand g347(n486, op1_i[1], op2_i[1]);
nand g348(product_o[1], n178, xenc101);
nand g349(n179, op2_i[1], op1_i[0]);
nand g350(n178, op2_i[0], op1_i[1]);
and g351(xenc0, n175, keyinput0);
or g352(xenc1, n443, keyinput1);
and g353(xenc2, n207, keyinput2);
and g354(xenc3, n470, keyinput3);
or g355(xenc4, n305, keyinput4);
or g356(xenc5, n312, keyinput5);
and g357(xenc6, n471, keyinput6);
or g358(xenc7, n423, keyinput7);
and g359(xenc8, n474, keyinput8);
and g360(xenc9, n379, keyinput9);
or g361(xenc10, n428, keyinput10);
and g362(xenc11, n451, keyinput11);
or g363(xenc12, n482, keyinput12);
or g364(xenc13, n410, keyinput13);
or g365(xenc14, n233, keyinput14);
and g366(xenc15, n402, keyinput15);
and g367(product_o[6], xenc16, keyinput16);
or g368(xenc17, n267, keyinput17);
or g369(product_o[10], xenc18, keyinput18);
and g370(xenc19, n357, keyinput19);
or g371(xenc20, n458, keyinput20);
or g372(xenc21, n468, keyinput21);
and g373(xenc22, n444, keyinput22);
or g374(xenc23, n367, keyinput23);
and g375(xenc24, n331, keyinput24);
and g376(xenc25, n243, keyinput25);
or g377(xenc26, n226, keyinput26);
and g378(xenc27, n480, keyinput27);
and g379(xenc28, n232, keyinput28);
and g380(xenc29, n419, keyinput29);
or g381(xenc30, n329, keyinput30);
and g382(xenc31, n344, keyinput31);
or g383(xenc32, n309, keyinput32);
or g384(xenc33, n347, keyinput33);
and g385(xenc34, n369, keyinput34);
and g386(xenc35, n144, keyinput35);
and g387(xenc36, n302, keyinput36);
and g388(xenc37, n368, keyinput37);
and g389(xenc38, n251, keyinput38);
and g390(xenc39, n194, keyinput39);
and g391(xenc40, n148, keyinput40);
or g392(product_o[7], xenc41, keyinput41);
and g393(xenc42, n236, keyinput42);
or g394(xenc43, n306, keyinput43);
and g395(xenc44, n418, keyinput44);
or g396(xenc45, n264, keyinput45);
and g397(xenc46, n403, keyinput46);
or g398(xenc47, n295, keyinput47);
or g399(xenc48, n449, keyinput48);
or g400(xenc49, n180, keyinput49);
or g401(xenc50, n384, keyinput50);
and g402(xenc51, n273, keyinput51);
and g403(xenc52, n422, keyinput52);
or g404(xenc53, n208, keyinput53);
or g405(xenc54, n364, keyinput54);
and g406(xenc55, n183, keyinput55);
or g407(xenc56, n326, keyinput56);
or g408(xenc57, n213, keyinput57);
and g409(xenc58, n206, keyinput58);
or g410(xenc59, n398, keyinput59);
or g411(xenc60, n465, keyinput60);
or g412(product_o[3], xenc61, keyinput61);
or g413(xenc62, n257, keyinput62);
and g414(product_o[2], xenc63, keyinput63);
and g415(xenc64, n397, keyinput64);
or g416(xenc65, n318, keyinput65);
and g417(xenc66, n231, keyinput66);
and g418(xenc67, n417, keyinput67);
or g419(xenc68, n427, keyinput68);
and g420(xenc69, n265, keyinput69);
or g421(xenc70, n307, keyinput70);
or g422(xenc71, n188, keyinput71);
or g423(xenc72, n254, keyinput72);
or g424(xenc73, n304, keyinput73);
or g425(xenc74, n200, keyinput74);
and g426(xenc75, n366, keyinput75);
or g427(xenc76, n242, keyinput76);
or g428(xenc77, n479, keyinput77);
or g429(xenc78, n247, keyinput78);
and g430(xenc79, n145, keyinput79);
and g431(xenc80, n212, keyinput80);
and g432(product_o[8], xenc81, keyinput81);
and g433(xenc82, n375, keyinput82);
and g434(xenc83, n420, keyinput83);
or g435(xenc84, n401, keyinput84);
or g436(xenc85, n313, keyinput85);
and g437(xenc86, n275, keyinput86);
or g438(xenc87, n485, keyinput87);
and g439(xenc88, n211, keyinput88);
or g440(xenc89, n230, keyinput89);
and g441(xenc90, n424, keyinput90);
or g442(xenc91, n291, keyinput91);
and g443(xenc92, n390, keyinput92);
and g444(xenc93, n395, keyinput93);
or g445(xenc94, n438, keyinput94);
or g446(xenc95, n256, keyinput95);
or g447(xenc96, n222, keyinput96);
and g448(xenc97, n340, keyinput97);
or g449(xenc98, n370, keyinput98);
or g450(product_o[11], xenc99, keyinput99);
and g451(xenc100, n198, keyinput100);
and g452(xenc101, n179, keyinput101);
and g453(xenc102, n314, keyinput102);
and g454(xenc103, n362, keyinput103);
and g455(xenc104, n260, keyinput104);
or g456(xenc105, n450, keyinput105);
and g457(xenc106, n282, keyinput106);
or g458(xenc107, n149, keyinput107);
and g459(xenc108, n322, keyinput108);
or g460(xenc109, n268, keyinput109);
or g461(xenc110, n350, keyinput110);
and g462(xenc111, n433, keyinput111);
or g463(xenc112, n388, keyinput112);
or g464(xenc113, n394, keyinput113);
and g465(xenc114, n164, keyinput114);
and g466(xenc115, n234, keyinput115);
and g467(xenc116, n315, keyinput116);
or g468(product_o[15], xenc117, keyinput117);
or g469(xenc118, n262, keyinput118);
or g470(xenc119, n162, keyinput119);
and g471(xenc120, n147, keyinput120);
and g472(xenc121, n219, keyinput121);
and g473(xenc122, n346, keyinput122);
and g474(xenc123, n440, keyinput123);
and g475(xenc124, n261, keyinput124);
and g476(xenc125, n203, keyinput125);
or g477(xenc126, n431, keyinput126);
or g478(product_o[5], xenc127, keyinput127);
endmodule
