module lower_part_or_ripple_carry_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  xor U95 ( result_o[9], n101, n102);
  xor U96 ( n102, add2_i[9], add1_i[9]);
  xor U97 ( result_o[8], add2_i[8], n103);
  xor U98 ( result_o[31], add2_i[31], n106);
  xor U100 ( result_o[30], add2_i[30], n110);
  xor U102 ( result_o[29], add2_i[29], n114);
  xor U104 ( result_o[28], add2_i[28], n118);
  xor U106 ( result_o[27], add2_i[27], n122);
  xor U108 ( result_o[26], add2_i[26], n126);
  xor U110 ( result_o[25], add2_i[25], n130);
  xor U111 ( n130, n131, add1_i[25]);
  xor U112 ( result_o[24], add2_i[24], n134);
  xor U114 ( result_o[23], add2_i[23], n138);
  xor U116 ( result_o[22], add2_i[22], n142);
  xor U118 ( result_o[21], add2_i[21], n146);
  xor U120 ( result_o[20], add2_i[20], n150);
  xor U122 ( result_o[19], add2_i[19], n154);
  xor U124 ( result_o[18], add2_i[18], n158);
  xor U126 ( result_o[17], add2_i[17], n162);
  xor U128 ( result_o[16], add2_i[16], n166);
  xor U130 ( result_o[15], add2_i[15], n170);
  xor U132 ( result_o[14], add2_i[14], n174);
  xor U134 ( result_o[13], add2_i[13], n178);
  xor U136 ( result_o[12], n182, add2_i[12]);
  xor U137 ( n182, n183, add1_i[12]);
  xor U138 ( result_o[11], n186, add2_i[11]);
  xor U139 ( n186, n187, add1_i[11]);
  xor U140 ( result_o[10], n190, add2_i[10]);
  xor U141 ( n190, n191, add1_i[10]);
  not U142 ( n199, add1_i[26]);
  not U143 ( n201, add1_i[24]);
  not U144 ( n198, add1_i[23]);
  xnor U145 ( n138, n139, n198);
  xnor U146 ( n126, n127, n199);
  not U147 ( n205, add1_i[22]);
  not U148 ( n200, add1_i[21]);
  xnor U149 ( n146, n147, n200);
  xnor U150 ( n134, n135, n201);
  not U151 ( n208, add1_i[20]);
  not U152 ( n203, add1_i[19]);
  not U153 ( n202, add1_i[29]);
  not U154 ( n204, add1_i[27]);
  xnor U155 ( n114, n115, n202);
  xnor U156 ( n154, n155, n203);
  xnor U157 ( n122, n123, n204);
  xnor U158 ( n142, n143, n205);
  not U159 ( n211, add1_i[18]);
  not U160 ( n206, add1_i[17]);
  not U161 ( n207, add1_i[28]);
  xnor U162 ( n162, n163, n206);
  xnor U163 ( n118, n119, n207);
  xnor U164 ( n150, n151, n208);
  not U165 ( n213, add1_i[31]);
  not U166 ( n209, add1_i[15]);
  not U167 ( n210, add1_i[30]);
  xnor U168 ( n170, n171, n209);
  xnor U169 ( n110, n111, n210);
  xnor U170 ( n158, n159, n211);
  not U171 ( n212, add1_i[16]);
  xnor U172 ( n166, n167, n212);
  xnor U173 ( n106, n107, n213);
  not U174 ( n214, add1_i[14]);
  not U175 ( n215, add1_i[13]);
  nand U176 ( n188, add1_i[10], n216);
  or U177 ( result_o[0], add1_i[0], add2_i[0]);
  or U178 ( result_o[1], add1_i[1], add2_i[1]);
  or U179 ( result_o[2], add1_i[2], add2_i[2]);
  or U180 ( result_o[3], add1_i[3], add2_i[3]);
  or U181 ( result_o[4], add1_i[4], add2_i[4]);
  or U182 ( result_o[5], add1_i[5], add2_i[5]);
  or U183 ( result_o[6], add1_i[6], add2_i[6]);
  nand U184 ( n184, add1_i[11], n187);
  xnor U185 ( n174, n175, n214);
  xnor U186 ( n178, n179, n215);
  or U187 ( result_o[7], add2_i[7], add1_i[7]);
  nand U188 ( n196, add1_i[8], add1_i[7], add2_i[7]);
  nand U189 ( n216, n192, n193);
  nand U190 ( n191, n193, n192);
  nand U191 ( n193, n194, add2_i[9]);
  nand U192 ( n180, n183, add1_i[12]);
  nand U193 ( n183, n185, n184);
  nand U194 ( n104, n107, add1_i[31]);
  nand U195 ( n107, n109, n108);
  nand U196 ( n197, add2_i[7], add1_i[7]);
  nand U197 ( n108, add1_i[30], n111);
  nand U198 ( n156, add1_i[18], n159);
  xnor U199 ( n103, n197, add1_i[8]);
  nand U200 ( n111, n112, n113);
  nand U201 ( n112, add1_i[29], n115);
  nand U202 ( n101, n195, n196);
  nand U203 ( n187, n188, n189);
  nand U204 ( n159, n160, n161);
  nand U205 ( n115, n116, n117);
  nand U206 ( n128, add1_i[25], n131);
  nand U207 ( n152, add1_i[19], n155);
  nand U208 ( n160, add1_i[17], n163);
  nand U209 ( n164, add1_i[16], n167);
  nand U210 ( n155, n156, n157);
  nand U211 ( n131, n132, n133);
  nand U212 ( n167, n168, n169);
  nand U213 ( n163, n164, n165);
  nand U214 ( n120, add1_i[27], n123);
  nand U215 ( n124, add1_i[26], n127);
  nand U216 ( n136, add1_i[23], n139);
  nand U217 ( n123, n124, n125);
  nand U218 ( n127, n128, n129);
  nand U219 ( n139, n140, n141);
  nand U220 ( n140, add1_i[22], n143);
  nand U221 ( n168, add1_i[15], n171);
  nand U222 ( n176, add1_i[13], n179);
  nand U223 ( n143, n144, n145);
  nand U224 ( n144, add1_i[21], n147);
  nand U225 ( n171, n172, n173);
  nand U226 ( n172, add1_i[14], n175);
  nand U227 ( n179, n180, n181);
  nand U228 ( n116, add1_i[28], n119);
  nand U229 ( n117, add2_i[28], n118);
  nand U230 ( n132, add1_i[24], n135);
  nand U231 ( n133, add2_i[24], n134);
  nand U232 ( n147, n148, n149);
  nand U233 ( n148, add1_i[20], n151);
  nand U234 ( n175, n176, n177);
  nand U235 ( n181, add2_i[12], n182);
  nand U236 ( result_o[32], n104, n105);
  nand U237 ( n105, add2_i[31], n106);
  nand U238 ( n119, n120, n121);
  nand U239 ( n129, add2_i[25], n130);
  nand U240 ( n135, n136, n137);
  nand U241 ( n145, add2_i[21], n146);
  nand U242 ( n151, n152, n153);
  nand U243 ( n157, add2_i[18], n158);
  nand U244 ( n169, add2_i[15], n170);
  nand U245 ( n192, add1_i[9], n101);
  or U246 ( n194, n101, add1_i[9]);
  nand U247 ( n195, n103, add2_i[8]);
  nand U248 ( n185, add2_i[11], n186);
  nand U249 ( n189, add2_i[10], n190);
  nand U250 ( n113, add2_i[29], n114);
  nand U251 ( n109, add2_i[30], n110);
  nand U252 ( n125, add2_i[26], n126);
  nand U253 ( n121, add2_i[27], n122);
  nand U254 ( n141, add2_i[22], n142);
  nand U255 ( n137, add2_i[23], n138);
  nand U256 ( n153, add2_i[19], n154);
  nand U257 ( n149, add2_i[20], n150);
  nand U258 ( n165, add2_i[16], n166);
  nand U259 ( n161, add2_i[17], n162);
  nand U260 ( n177, add2_i[13], n178);
  nand U261 ( n173, add2_i[14], n174);
endmodule
