module lower_part_or_ripple_carry_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83;

  xor U50 ( result_o[9], add2_i[9], n36);
  xor U51 ( result_o[8], add2_i[8], n37);
  xor U52 ( result_o[7], add2_i[7], n38);
  xor U53 ( result_o[6], add2_i[6], n39);
  xor U54 ( result_o[5], add2_i[5], n40);
  xor U55 ( result_o[4], add2_i[4], n41);
  xor U56 ( result_o[15], add2_i[15], n44);
  xor U57 ( n44, n45, add1_i[15]);
  xor U58 ( result_o[14], add2_i[14], n48);
  xor U59 ( n48, n49, add1_i[14]);
  xor U60 ( result_o[13], add2_i[13], n52);
  xor U61 ( n52, n53, add1_i[13]);
  xor U62 ( result_o[12], add2_i[12], n56);
  xor U63 ( n56, n57, add1_i[12]);
  xor U64 ( result_o[11], add2_i[11], n60);
  xor U65 ( n60, n61, add1_i[11]);
  xor U66 ( result_o[10], add2_i[10], n64);
  xor U67 ( n64, n65, add1_i[10]);
  xor U68 ( n36, n68, add1_i[9]);
  xor U69 ( n37, n71, add1_i[8]);
  xor U70 ( n38, n74, add1_i[7]);
  xor U71 ( n39, n77, add1_i[6]);
  xor U72 ( n40, n80, add1_i[5]);
  xnor U73 ( n41, n83, add1_i[4]);
  nand U74 ( n83, add2_i[3], add1_i[3]);
  nand U75 ( n77, n78, n79);
  nand U76 ( n78, add1_i[5], n80);
  nand U77 ( n79, add2_i[5], n40);
  nand U78 ( n74, n75, n76);
  nand U79 ( n75, add1_i[6], n77);
  nand U80 ( n76, add2_i[6], n39);
  nand U81 ( n53, n54, n55);
  nand U82 ( n54, add1_i[12], n57);
  nand U83 ( n55, add2_i[12], n56);
  nand U84 ( n49, n50, n51);
  nand U85 ( n50, add1_i[13], n53);
  nand U86 ( n51, add2_i[13], n52);
  nand U87 ( n45, n46, n47);
  nand U88 ( n46, add1_i[14], n49);
  nand U89 ( n47, add2_i[14], n48);
  nand U90 ( n80, n81, n82);
  nand U91 ( n82, add1_i[4], add1_i[3], add2_i[3]);
  nand U92 ( n81, add2_i[4], n41);
  nand U93 ( n71, n72, n73);
  nand U94 ( n72, add1_i[7], n74);
  nand U95 ( n73, add2_i[7], n38);
  nand U96 ( n68, n69, n70);
  nand U97 ( n69, add1_i[8], n71);
  nand U98 ( n70, add2_i[8], n37);
  nand U99 ( n65, n66, n67);
  nand U100 ( n66, add1_i[9], n68);
  nand U101 ( n67, add2_i[9], n36);
  nand U102 ( n61, n62, n63);
  nand U103 ( n62, add1_i[10], n65);
  nand U104 ( n63, add2_i[10], n64);
  nand U105 ( n57, n58, n59);
  nand U106 ( n58, add1_i[11], n61);
  nand U107 ( n59, add2_i[11], n60);
  nand U108 ( result_o[16], n42, n43);
  nand U109 ( n42, add1_i[15], n45);
  nand U110 ( n43, add2_i[15], n44);
  or U111 ( result_o[0], add1_i[0], add2_i[0]);
  or U112 ( result_o[1], add1_i[1], add2_i[1]);
  or U113 ( result_o[2], add1_i[2], add2_i[2]);
  or U114 ( result_o[3], add2_i[3], add1_i[3]);
endmodule
