library verilog;
use verilog.vl_types.all;
entity equal_segmentation_adder32_tb is
end equal_segmentation_adder32_tb;
