module equal_segmentation_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;

  xor U36 ( result_o[9], add2_i[9], n28);
  xor U37 ( result_o[8], add2_i[8], add1_i[8]);
  xor U38 ( result_o[7], n29, n30);
  xor U39 ( n30, add2_i[7], add1_i[7]);
  xor U40 ( result_o[6], add2_i[6], n33);
  xor U41 ( n33, n34, add1_i[6]);
  xor U42 ( result_o[5], add2_i[5], n37);
  xor U43 ( result_o[4], add2_i[4], add1_i[4]);
  xor U44 ( result_o[3], n39, n40);
  xor U45 ( n40, add2_i[3], add1_i[3]);
  xor U46 ( result_o[2], add2_i[2], n43);
  xor U47 ( n43, n44, add1_i[2]);
  xor U48 ( result_o[1], add2_i[1], n47);
  xor U49 ( result_o[15], add2_i[15], n51);
  xor U50 ( n51, n52, add1_i[15]);
  xor U51 ( result_o[14], add2_i[14], n55);
  xor U52 ( n55, n56, add1_i[14]);
  xor U53 ( result_o[13], add2_i[13], n59);
  xor U54 ( result_o[12], add2_i[12], add1_i[12]);
  xor U55 ( result_o[11], n61, n62);
  xor U56 ( n62, add2_i[11], add1_i[11]);
  xor U57 ( result_o[10], add2_i[10], n65);
  xor U58 ( n65, n66, add1_i[10]);
  xor U59 ( result_o[0], add2_i[0], add1_i[0]);
  xnor U60 ( n59, n60, add1_i[13]);
  nand U61 ( n60, add2_i[12], add1_i[12]);
  xnor U62 ( n47, n48, add1_i[1]);
  nand U63 ( n48, add2_i[0], add1_i[0]);
  xnor U64 ( n37, n38, add1_i[5]);
  nand U65 ( n38, add2_i[4], add1_i[4]);
  xnor U66 ( n28, n69, add1_i[9]);
  nand U67 ( n69, add2_i[8], add1_i[8]);
  nand U68 ( n39, n41, n42);
  nand U69 ( n41, add1_i[2], n44);
  nand U70 ( n29, n31, n32);
  nand U71 ( n31, add1_i[6], n34);
  nand U72 ( n61, n63, n64);
  nand U73 ( n63, add1_i[10], n66);
  nand U74 ( n52, n53, n54);
  nand U75 ( n53, add1_i[14], n56);
  nand U76 ( n54, add2_i[14], n55);
  nand U77 ( n42, add2_i[2], n43);
  nand U78 ( n32, add2_i[6], n33);
  nand U79 ( n64, add2_i[10], n65);
  nand U80 ( n56, n57, n58);
  nand U81 ( n58, add1_i[13], add1_i[12], add2_i[12]);
  nand U82 ( n57, add2_i[13], n59);
  nand U83 ( n44, n45, n46);
  nand U84 ( n46, add1_i[1], add1_i[0], add2_i[0]);
  nand U85 ( n45, add2_i[1], n47);
  nand U86 ( n34, n35, n36);
  nand U87 ( n36, add1_i[5], add1_i[4], add2_i[4]);
  nand U88 ( n35, add2_i[5], n37);
  nand U89 ( n66, n67, n68);
  nand U90 ( n68, add2_i[8], add1_i[8], add1_i[9]);
  nand U91 ( n67, add2_i[9], n28);
  nand U92 ( result_o[16], n49, n50);
  nand U93 ( n49, add1_i[15], n52);
  nand U94 ( n50, add2_i[15], n51);
endmodule
