library verilog;
use verilog.vl_types.all;
entity lower_part_or_carry_lookahead_adder16_tb is
end lower_part_or_carry_lookahead_adder16_tb;
