module underdesigned_multiplier8 ( op1_i, op2_i, product_o );
  input [7:0] op1_i, op2_i;
  output [15:0] product_o;
  wire   n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n166, n167, n169, n170, n171, n172, n173, n174, n175, n177, n178,
         n179, n180, n181, n182, n183, n184, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486;

  xor U310 ( product_o[9], n158, n159);
  xor U311 ( product_o[8], n160, n161);
  xor U312 ( n160, n162, n163);
  xor U314 ( product_o[5], n171, n170);
  xor U315 ( product_o[3], n174, n175);
  xor U318 ( n183, n186, n187);
  xor U321 ( n232, n236, n208);
  xor U323 ( n221, n229, n230);
  xor U324 ( n229, n234, n235);
  xor U326 ( n272, n274, n275);
  xor U327 ( n268, n298, n261);
  xor U328 ( n169, n320, n319);
  xor U329 ( n320, n332, n333);
  xor U330 ( n170, n327, n331);
  xor U331 ( n331, n334, n335);
  xor U332 ( n329, n336, n337);
  xor U333 ( n338, n340, n341);
  xor U334 ( n343, n346, n347);
  xor U335 ( n332, n350, n351);
  xor U336 ( n347, n352, n353);
  xor U337 ( n335, n354, n355);
  xor U338 ( n354, n356, n357);
  xor U339 ( n352, n380, n381);
  xor U340 ( n381, n382, n383);
  xor U341 ( n353, n378, n379);
  xor U342 ( n159, n314, n313);
  xor U343 ( n368, n396, n391);
  xor U344 ( n396, n392, n389);
  xor U345 ( n385, n415, n416);
  xor U346 ( n386, n417, n418);
  xor U347 ( n312, n289, n288);
  xor U348 ( n309, n303, n422);
  xor U349 ( n455, n456, n457);
  xor U351 ( n417, n462, n435);
  xor U352 ( n420, n470, n441);
  nand U353 ( n215, n243, n244);
  nand U354 ( n243, n247, n245);
  nand U355 ( n244, n245, n246);
  and U356 ( n278, n159, n158);
  nand U357 ( n246, n276, n277);
  nand U358 ( n276, n280, n279);
  nand U359 ( n277, n278, n279);
  xnor U360 ( product_o[10], n478, n279);
  nor U361 ( n478, n278, n280);
  xnor U362 ( product_o[11], n479, n245);
  nor U363 ( n479, n246, n247);
  nor U364 ( n279, n247, n282);
  and U365 ( n282, n283, n284);
  nor U366 ( n247, n284, n283);
  nand U367 ( n316, n353, n352, n149);
  not U368 ( n149, n374);
  nand U369 ( n167, n319, n320);
  xnor U370 ( product_o[13], n480, n194);
  nor U371 ( n480, n195, n143);
  nand U372 ( n162, n164, n318);
  nand U373 ( n318, n166, n167);
  nand U374 ( n158, n315, n316);
  nand U375 ( n315, n163, n317);
  nand U376 ( n317, n161, n162);
  nand U377 ( n184, n192, n193);
  nand U378 ( n192, n143, n194);
  nand U379 ( n193, n194, n195);
  and U380 ( n163, n316, n372);
  nand U381 ( n372, n373, n374);
  nand U382 ( n373, n353, n352);
  nor U383 ( n245, n216, n249);
  and U384 ( n249, n250, n251);
  nor U385 ( n216, n251, n250);
  xnor U386 ( n250, n222, n221);
  nor U387 ( n280, n313, n314);
  xor U388 ( product_o[7], n164, n481);
  nand U389 ( n481, n166, n167);
  xnor U390 ( n418, n419, n420);
  xnor U391 ( n333, n348, n349);
  nand U392 ( n348, n335, n334);
  xnor U393 ( n164, n342, n343);
  nand U394 ( n342, n332, n333);
  xnor U395 ( n286, n272, n273);
  nand U396 ( n166, n170, n169, n171);
  nand U397 ( n251, n289, n288, n148);
  not U398 ( n148, n286);
  nand U399 ( n313, n379, n378, n377);
  nand U400 ( n419, n447, n448);
  or U401 ( n447, n382, n383);
  nand U402 ( n448, n380, n449);
  nand U403 ( n449, n383, n382);
  nand U404 ( n294, n444, n445);
  or U405 ( n444, n420, n417);
  nand U406 ( n445, n446, n419);
  nand U407 ( n446, n417, n420);
  nand U408 ( n275, n291, n292);
  nand U409 ( n291, n295, n296);
  nand U410 ( n292, n293, n294);
  or U411 ( n293, n295, n296);
  nand U412 ( n283, n251, n285);
  nand U413 ( n285, n286, n287);
  nand U414 ( n287, n288, n289);
  and U415 ( n161, n344, n345);
  nand U416 ( n344, n346, n347);
  nand U417 ( n345, n332, n333, n343);
  nand U418 ( n195, n212, n213);
  nand U419 ( n212, n216, n214);
  nand U420 ( n213, n214, n215);
  nand U421 ( n374, n313, n375);
  nand U422 ( n375, n376, n150);
  nand U423 ( n376, n378, n379);
  not U424 ( n150, n377);
  xnor U425 ( n289, n431, n295);
  xnor U426 ( n431, n294, n296);
  nor U427 ( n194, n182, n197);
  and U428 ( n197, n198, n199);
  nor U429 ( n182, n199, n198);
  xnor U430 ( n314, n312, n311);
  nand U431 ( n200, n229, n230, n145);
  not U432 ( n145, n228);
  nand U433 ( n191, n235, n234, n147);
  not U434 ( n147, n232);
  nand U435 ( n222, n270, n271);
  nand U436 ( n270, n274, n275);
  nand U437 ( n271, n272, n273);
  xnor U438 ( product_o[6], n482, n169);
  nand U439 ( n482, n170, n171);
  nand U440 ( n225, n200, n226);
  nand U441 ( n226, n227, n228);
  nand U442 ( n227, n229, n230);
  nand U443 ( n284, n311, n312);
  xnor U444 ( product_o[12], n483, n214);
  nor U445 ( n483, n215, n216);
  nand U446 ( n228, n191, n231);
  nand U447 ( n231, n232, n233);
  nand U448 ( n233, n234, n235);
  not U449 ( n143, n211);
  and U450 ( n319, n327, n331);
  and U451 ( n198, n200, n201);
  and U452 ( n346, n349, n334, n335);
  xnor U453 ( n470, n443, n442);
  xnor U454 ( n422, n304, n302);
  nor U455 ( n402, n153, n409, n155);
  nor U456 ( n452, n151, n157, n460);
  nor U457 ( n304, n154, n152, n425);
  nor U458 ( n311, n386, n385);
  xnor U459 ( n349, n368, n369);
  xnor U460 ( n369, n370, n371);
  xnor U461 ( n383, n454, n455);
  xnor U462 ( n337, n409, n414);
  nor U463 ( n414, n153, n155);
  nor U464 ( n377, n311, n384);
  and U465 ( n384, n385, n386);
  xnor U466 ( n274, n297, n268);
  xnor U467 ( n297, n267, n269);
  nor U468 ( n458, n155, n152);
  xnor U469 ( n380, n450, n451);
  xnor U470 ( n451, n452, n453);
  xnor U471 ( n355, n401, n406);
  xnor U472 ( n406, n402, n400);
  nand U473 ( n379, n393, n394);
  or U474 ( n393, n370, n371);
  nand U475 ( n394, n368, n395);
  nand U476 ( n395, n371, n370);
  and U477 ( n371, n403, n404);
  or U478 ( n403, n356, n357);
  nand U479 ( n404, n355, n405);
  nand U480 ( n405, n357, n356);
  nand U481 ( n267, n305, n306);
  or U482 ( n305, n310, n309);
  nand U483 ( n306, n307, n308);
  nand U484 ( n307, n309, n310);
  xnor U485 ( product_o[14], n484, n183);
  nor U486 ( n484, n184, n182);
  nand U487 ( n441, n471, n472);
  or U488 ( n471, n456, n454);
  nand U489 ( n472, n473, n457);
  nand U490 ( n473, n454, n456);
  and U491 ( n391, n397, n398);
  nand U492 ( n397, n402, n401);
  nand U493 ( n398, n399, n400);
  or U494 ( n399, n401, n402);
  nand U495 ( product_o[15], n180, n181);
  nand U496 ( n181, n182, n183);
  nand U497 ( n180, n183, n184);
  xnor U498 ( n298, n263, n262);
  xnor U499 ( n462, n437, n436);
  nor U500 ( n242, n151, n155, n255);
  nor U501 ( n325, n153, n156, n321);
  xnor U502 ( n236, n210, n209);
  xnor U503 ( n175, n323, n324);
  xnor U504 ( n324, n325, n326);
  xnor U505 ( n230, n241, n252);
  xnor U506 ( n252, n242, n240);
  xnor U507 ( n288, n421, n309);
  xnor U508 ( n421, n310, n308);
  xnor U509 ( n273, n255, n290);
  nor U510 ( n290, n155, n151);
  nor U511 ( n327, n330, n329);
  nor U512 ( n172, n327, n328);
  and U513 ( n328, n329, n330);
  xnor U514 ( n177, n321, n322);
  nor U515 ( n322, n156, n153);
  xnor U516 ( n416, n425, n430);
  nor U517 ( n430, n152, n154);
  nand U518 ( n211, n221, n222, n144);
  not U519 ( n144, n220);
  xnor U520 ( n330, n338, n339);
  xnor U521 ( n199, n190, n189);
  xnor U522 ( n351, n460, n461);
  nor U523 ( n461, n157, n151);
  nand U524 ( n296, n438, n439);
  or U525 ( n438, n443, n442);
  nand U526 ( n439, n440, n441);
  nand U527 ( n440, n442, n443);
  nand U528 ( n295, n432, n433);
  or U529 ( n432, n437, n436);
  nand U530 ( n433, n434, n435);
  nand U531 ( n434, n436, n437);
  nand U532 ( n334, n358, n359);
  or U533 ( n358, n340, n339);
  nand U534 ( n359, n341, n360);
  nand U535 ( n360, n339, n340);
  nand U536 ( n235, n258, n259);
  or U537 ( n258, n262, n263);
  nand U538 ( n259, n260, n261);
  nand U539 ( n260, n262, n263);
  and U540 ( n339, n361, n362);
  nand U541 ( n361, n325, n323);
  nand U542 ( n362, n363, n326);
  or U543 ( n363, n323, n325);
  nand U544 ( n378, n387, n388);
  or U545 ( n387, n392, n391);
  nand U546 ( n388, n389, n390);
  nand U547 ( n390, n391, n392);
  nand U548 ( n234, n264, n265);
  or U549 ( n264, n269, n268);
  nand U550 ( n265, n266, n267);
  nand U551 ( n266, n268, n269);
  and U552 ( n214, n211, n218);
  nand U553 ( n218, n219, n220);
  nand U554 ( n219, n221, n222);
  nor U555 ( n188, n189, n190);
  nand U556 ( n190, n204, n191);
  nand U557 ( n204, n205, n206);
  or U558 ( n205, n210, n209);
  nand U559 ( n206, n207, n208);
  nand U560 ( n382, n351, n350);
  nand U561 ( n435, n463, n464);
  nand U562 ( n463, n452, n450);
  nand U563 ( n464, n465, n453);
  or U564 ( n465, n450, n452);
  nand U565 ( n261, n299, n300);
  nand U566 ( n299, n304, n303);
  nand U567 ( n300, n301, n302);
  or U568 ( n301, n303, n304);
  nand U569 ( n208, n237, n238);
  nand U570 ( n237, n242, n241);
  nand U571 ( n238, n239, n240);
  or U572 ( n239, n241, n242);
  and U573 ( n171, n172, n175, n174);
  or U574 ( n201, n151, n154, n225);
  nand U575 ( n207, n209, n210);
  xnor U576 ( product_o[4], n172, n173);
  nand U577 ( n173, n174, n175);
  nor U578 ( product_o[0], n153, n157);
  not U579 ( n153, op1_i[0]);
  not U580 ( n155, op2_i[4]);
  nand U581 ( n356, op1_i[4], n337, op2_i[0]);
  nand U582 ( n456, op1_i[4], op2_i[2], n458);
  nand U583 ( n401, n410, n411);
  nand U584 ( n410, op2_i[4], op1_i[1]);
  nand U585 ( n411, op1_i[0], op2_i[5]);
  not U586 ( n152, op1_i[2]);
  nand U587 ( n400, n407, n408);
  nand U588 ( n407, op2_i[2], op1_i[3]);
  nand U589 ( n408, op1_i[2], op2_i[3]);
  nand U590 ( n409, op2_i[2], op1_i[2]);
  nand U591 ( n460, op2_i[6], op1_i[0]);
  nand U592 ( n425, op1_i[4], op2_i[4]);
  nand U593 ( n186, op1_i[7], op2_i[7]);
  nor U594 ( n187, n146, n188);
  not U595 ( n146, n191);
  xnor U596 ( n350, n458, n485);
  nand U597 ( n485, op2_i[2], op1_i[4]);
  nand U598 ( n415, op1_i[6], op2_i[2]);
  nand U599 ( n336, op2_i[0], op1_i[4]);
  not U600 ( n151, op1_i[6]);
  nand U601 ( n310, op2_i[2], n416, op1_i[6]);
  nand U602 ( n269, op1_i[7], op2_i[3]);
  nand U603 ( n443, op2_i[5], op1_i[3]);
  nand U604 ( n437, op2_i[7], op1_i[1]);
  nand U605 ( n370, op2_i[1], op1_i[5]);
  nand U606 ( n210, op2_i[7], op1_i[5]);
  nand U607 ( n323, n366, n367);
  nand U608 ( n366, op2_i[2], op1_i[1]);
  nand U609 ( n367, op1_i[0], op2_i[3]);
  nand U610 ( n450, n468, n469);
  nand U611 ( n468, op2_i[6], op1_i[1]);
  nand U612 ( n469, op2_i[7], op1_i[0]);
  nand U613 ( n241, n256, n257);
  nand U614 ( n256, op2_i[6], op1_i[5]);
  nand U615 ( n257, op2_i[7], op1_i[4]);
  nand U616 ( n262, op2_i[7], op1_i[3]);
  nand U617 ( n263, op1_i[5], op2_i[5]);
  nand U618 ( n442, op1_i[5], op2_i[3]);
  nand U619 ( n436, op1_i[7], op2_i[1]);
  nand U620 ( n209, op1_i[7], op2_i[5]);
  not U621 ( n154, op2_i[6]);
  not U622 ( n157, op2_i[0]);
  and U623 ( n454, n476, n477);
  nand U624 ( n476, op2_i[4], op1_i[3]);
  nand U625 ( n477, op1_i[2], op2_i[5]);
  nand U626 ( n453, n466, n467);
  nand U627 ( n466, op1_i[7], op2_i[0]);
  nand U628 ( n467, op1_i[6], op2_i[1]);
  nand U629 ( n326, n364, n365);
  nand U630 ( n364, op2_i[0], op1_i[3]);
  nand U631 ( n365, op2_i[1], op1_i[2]);
  nand U632 ( n308, n428, n429);
  nand U633 ( n428, op1_i[7], op2_i[2]);
  nand U634 ( n429, op1_i[6], op2_i[3]);
  nand U635 ( n302, n423, n424);
  nand U636 ( n423, op2_i[6], op1_i[3]);
  nand U637 ( n424, op2_i[7], op1_i[2]);
  nand U638 ( n240, n253, n254);
  nand U639 ( n253, op1_i[7], op2_i[4]);
  nand U640 ( n254, op1_i[6], op2_i[5]);
  nand U641 ( n303, n426, n427);
  nand U642 ( n426, op1_i[5], op2_i[4]);
  nand U643 ( n427, op1_i[4], op2_i[5]);
  nand U644 ( n340, op1_i[1], op2_i[3]);
  nand U645 ( n392, op2_i[5], op1_i[1]);
  nand U646 ( n321, op2_i[0], op1_i[2]);
  nand U647 ( n255, op2_i[6], op1_i[4]);
  and U648 ( n357, n412, n413);
  nand U649 ( n412, op2_i[0], op1_i[5]);
  nand U650 ( n413, op1_i[4], op2_i[1]);
  nand U651 ( n220, n201, n223);
  nand U652 ( n223, n224, n225);
  nand U653 ( n224, op1_i[6], op2_i[6]);
  and U654 ( n174, op1_i[1], n177, op2_i[1]);
  and U655 ( n389, op2_i[3], op1_i[3]);
  and U656 ( n341, op2_i[1], op1_i[3]);
  not U657 ( n156, op2_i[2]);
  nand U658 ( n457, n474, n475);
  nand U659 ( n474, op1_i[5], op2_i[2]);
  nand U660 ( n475, op1_i[4], op2_i[3]);
  and U661 ( n189, n202, n203);
  nand U662 ( n202, op1_i[7], op2_i[6]);
  nand U663 ( n203, op2_i[7], op1_i[6]);
  xnor U664 ( product_o[2], n486, n177);
  nand U665 ( n486, op1_i[1], op2_i[1]);
  nand U666 ( product_o[1], n178, n179);
  nand U667 ( n179, op2_i[1], op1_i[0]);
  nand U668 ( n178, op2_i[0], op1_i[1]);
endmodule
