// Verilog File 
module ripple_carry_adder32_xor_enc64.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,result_o[0],
result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],result_o[7],result_o[8],result_o[9],result_o[10],
result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],result_o[17],result_o[18],result_o[19],result_o[20],
result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],result_o[27],result_o[28],result_o[29],result_o[30],
result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n886, xenc16, n812, n816, n817, xenc10, xenc42, xenc57, n820, 
n837, xenc48, xenc31, n846, xenc18, n857, xenc38, n859, xenc8, n863, 
n864, n867, xenc63, n871, xenc23, n875, xenc26, xenc32, xenc2, n887, 
xenc56, xenc59, n894, xenc19, n907, n912, n913, xenc41, xenc22, n926, 
xenc35, n927, xenc53, n960, n796, n992, n841, n1002, n915, n1001, 
n911, n836, n998, n995, n931, n977, xenc28, n959, n958, n957, 
n965, xenc36, n996, n800, n900, n901, n893, n966, n974, n928, 
xenc15, n988, n948, n985, n967, n1000, n865, n902, n969, n976, 
n830, n827, n937, xenc51, n938, xenc21, n921, n872, n855, n968, 
xenc58, n980, n840, n983, n818, n904, n903, n799, n896, n881, 
n880, n823, xenc40, n849, xenc61, n848, n1003, n970, n897, xenc30, 
n910, n971, n815, n936, n972, n973, xenc5, n925, xenc46, n860, 
n975, n941, xenc7, n892, n978, n890, n979, n990, n991, n981, 
n982, n986, n984, xenc25, n987, n918, n989, xenc13, xenc44, n916, 
n845, n847, n993, n933, n801, xenc1, n994, n831, n997, n999, 
n862, xenc37, n954, n1005, n1004, n930, n876, n1006, n1007, xenc33, 
n884, xenc49, n1012, n1011, n833, n834, n835, n851, n850, n852, 
n798, n853, n951, xenc62, xenc14, xenc45, n1008, n1009, n832, n802, 
xenc54, n939, n944, n940, xenc29, n945, n803, n898, n917, n1010, 
n814, xenc47, xenc52, n797, n947, n943, n888, n889, n885, xenc34, 
n879, n924, n923, n922, xenc0, n861, n825, n826, n824, xenc43, 
n956, n914, n955, n952, n873, xenc55, n919, xenc6, xenc60, n963, 
n962, n877, xenc3, n821, n866, n810, n932, n946, n839, xenc4, 
n869, n868, n905, n953, n819, n828, xenc20, n891, xenc17, xenc50, 
n935, n811, n934, n858, n856, n854, xenc27, n878, n929, n809, 
xenc24, n822, n808, n883, n882, n906, xenc12, n961, xenc39, n895, 
n870, n874, n909, n920, xenc9, xenc11, n942;

or g0(n886, add2_i[0], add1_i[0]);
xor g1(result_o[8], xenc16, n812);
xor g2(result_o[6], add2_i[6], n816);
xor g3(result_o[5], add2_i[5], n817);
xor g4(xenc57, xenc10, xenc42);
xor g5(n820, add2_i[3], add1_i[3]);
xor g6(xenc48, n837, add2_i[2]);
xor g7(result_o[28], add2_i[28], xenc31);
xor g8(result_o[27], add2_i[27], n846);
xor g9(xenc38, xenc18, n857);
xor g10(xenc8, n859, add2_i[25]);
xor g11(result_o[24], n863, n864);
xor g12(n864, add2_i[24], add1_i[24]);
xor g13(xenc63, add2_i[23], n867);
xor g14(xenc23, add2_i[22], n871);
xor g15(xenc26, add2_i[21], n875);
xor g16(xenc2, n886, xenc32);
xor g17(n887, add2_i[1], add1_i[1]);
xor g18(xenc59, xenc56, add2_i[19]);
xor g19(result_o[18], n894, xenc19);
xor g20(result_o[15], add2_i[15], n907);
xor g21(result_o[14], n912, n913);
xor g22(n913, add2_i[14], add1_i[14]);
xor g23(xenc22, xenc41, add2_i[12]);
xor g24(result_o[11], n926, xenc35);
xor g25(n927, add2_i[11], add1_i[11]);
xor g26(result_o[10], xenc53, add2_i[10]);
xor g27(n837, n960, add1_i[2]);
nand g28(n841, n796, n992);
nand g29(n911, n1002, n915, n1001);
nand g30(n995, n836, add2_i[28], add1_i[29], n998);
xor g31(n977, n931, add1_i[10]);
nand g32(n957, xenc28, n959, n958);
not g33(n965, add1_i[3]);
nand g34(n996, xenc36, add1_i[28], add1_i[29]);
nand g35(n893, n800, n900, n901);
nor g36(n974, n966, add1_i[11]);
not g37(n966, n928);
and g38(n985, xenc15, n988, n948);
nor g39(n1000, n967, add1_i[24]);
not g40(n967, n865);
nand g41(n969, n902, add2_i[16], add1_i[17]);
nand g42(n827, n976, n995, n996, n830);
nand g43(n938, n937, xenc51, add2_i[6]);
xor g44(n921, xenc21, add1_i[12]);
xor g45(n871, n872, add1_i[22]);
xor g46(n859, n855, add1_i[25]);
nor g47(n840, n968, xenc58, n980);
not g48(n968, n983);
xnor g49(result_o[0], add2_i[0], add1_i[0]);
xor g50(result_o[4], add2_i[4], n818);
xnor g51(n903, n904, add1_i[16]);
and g52(n896, add2_i[17], n893, n799);
xnor g53(n880, n881, add1_i[20]);
xor g54(xenc40, n823, add2_i[31]);
and g55(n848, n849, xenc61);
not g56(n1003, add1_i[4]);
nand g57(n897, n969, n970);
or g58(n970, n800, n901);
nand g59(n971, xenc30, n910);
nand g60(n972, n815, n936);
nand g61(n973, n977, add2_i[10]);
nand g62(n925, n973, xenc5);
nand g63(n975, xenc46, n860);
not g64(n976, add1_i[30]);
and g65(n815, n941, xenc7);
and g66(n816, xenc51, n937);
nand g67(n890, n892, n978);
nor g68(n978, n897, add1_i[18]);
and g69(n979, n817, n988);
nor g70(n998, n980, xenc58);
and g71(n980, add1_i[28], n990);
and g72(n981, n991, add1_i[28]);
or g73(n982, n991, add1_i[28], n990);
or g74(n983, n991, add1_i[28], n990);
or g75(n836, n991, add1_i[28], n990);
nor g76(n984, n979, n986);
nor g77(n937, n985, n986);
nor g78(n986, xenc25, xenc15);
not g79(n987, add1_i[6]);
and g80(n988, add2_i[5], add1_i[6]);
or g81(n989, n918, add1_i[13]);
nor g82(n990, n992, xenc13);
nor g83(n991, xenc44, n848);
or g84(n916, n918, add1_i[13]);
nor g85(n845, xenc44, n848);
nand g86(n992, add2_i[27], n847);
nand g87(n993, xenc30, n910);
nand g88(n994, n933, n801, xenc1);
and g89(n831, n995, n996);
not g90(n997, add1_i[29]);
nand g91(n999, n867, add2_i[23]);
nand g92(n862, n999, n1000);
nand g93(n1001, xenc37, add2_i[13]);
not g94(n1002, add1_i[14]);
xnor g95(n818, n954, n1003);
not g96(n1005, add1_i[21]);
not g97(n1004, add1_i[10]);
xnor g98(n930, n931, n1004);
xnor g99(n875, n876, n1005);
not g100(n1006, add1_i[19]);
not g101(n1007, add1_i[31]);
xnor g102(n884, xenc33, n1006);
xnor g103(n823, xenc49, n1007);
not g104(n1012, add1_i[15]);
not g105(n1011, add1_i[23]);
nand g106(n830, n833, add2_i[29]);
nand g107(n833, n834, n997, n835);
nand g108(n850, add2_i[26], n851);
nand g109(n851, n852, n798, n853);
not g110(n801, add1_i[9]);
xnor g111(n857, add2_i[26], n798);
or g112(n948, n951, add1_i[5]);
xor g113(xenc45, xenc62, xenc14);
xor g114(n1008, add1_i[30], add2_i[30]);
xor g115(result_o[29], n1009, n832);
xor g116(n1009, add1_i[29], add2_i[29]);
nand g117(n834, add1_i[28], xenc36);
not g118(n802, add1_i[8]);
xnor g119(xenc54, add2_i[20], n880);
nand g120(n933, add2_i[8], n939);
nand g121(n940, add2_i[7], n944);
nand g122(n852, add2_i[25], xenc29);
nand g123(n945, add2_i[6], xenc51);
not g124(n803, add1_i[7]);
xnor g125(n894, add1_i[18], add2_i[18]);
xnor g126(result_o[17], add2_i[17], n898);
xnor g127(result_o[13], add2_i[13], n917);
xnor g128(result_o[16], add2_i[16], n903);
not g129(n800, add1_i[17]);
xnor g130(n812, add2_i[8], n802);
not g131(n798, add1_i[26]);
xnor g132(result_o[7], add2_i[7], n1010);
nand g133(n1010, n814, n815);
xnor g134(xenc52, add2_i[9], xenc47);
not g135(n797, add1_i[27]);
nand g136(n943, xenc15, xenc25, n947);
nand g137(n885, n888, n889);
xnor g138(n867, xenc34, n1011);
xnor g139(n907, n993, n1012);
or g140(n902, n904, add1_i[16]);
or g141(n879, n881, add1_i[20]);
nand g142(n917, n915, xenc37);
nand g143(n910, n911, add2_i[14]);
nand g144(n924, n925, add2_i[11]);
nand g145(n922, n924, n923);
nand g146(n855, xenc46, n860);
nand g147(n861, add2_i[24], xenc0);
nand g148(n947, n948, add2_i[5]);
nand g149(n824, n825, n826);
nand g150(n956, xenc43, add2_i[3]);
nand g151(n914, n916, add2_i[13]);
and g152(n846, n796, n847);
nand g153(n826, n827, add2_i[30]);
and g154(n817, xenc15, n948);
nand g155(n958, add1_i[2], n960);
nand g156(n954, n956, n955);
nand g157(n952, add1_i[4], n954);
nand g158(n847, n848, xenc44);
nand g159(n873, add1_i[21], n876);
nand g160(n889, xenc55, add2_i[18]);
nand g161(n919, add1_i[12], xenc21);
nand g162(n912, n914, n915);
nand g163(n900, n902, add2_i[16]);
nand g164(n960, xenc6, xenc60);
nand g165(n962, n963, add2_i[1]);
nand g166(n876, n877, xenc3);
nand g167(n877, n879, add2_i[20]);
nand g168(n821, add1_i[31], xenc49);
nand g169(n863, n865, n866);
nand g170(n865, xenc34, add1_i[23]);
nand g171(n928, n931, add1_i[10]);
nand g172(n931, n810, n932);
nand g173(n939, n940, n802, n815);
nand g174(n946, add1_i[5], n951);
nand g175(n832, n834, n839);
nand g176(n868, xenc4, n869);
nand g177(n869, n872, add1_i[22]);
nand g178(n905, n971, add1_i[15]);
nand g179(n915, add1_i[13], n918);
nand g180(n951, n953, n952);
nand g181(n819, n959, n958);
nand g182(n828, n831, n830);
nand g183(n839, add2_i[28], xenc31);
nand g184(n849, add1_i[26], xenc18);
nand g185(n888, add1_i[18], xenc20);
nand g186(n891, n892, n799);
nand g187(n918, xenc17, xenc50);
nand g188(n810, n935, add1_i[9]);
nand g189(n934, add1_i[8], n811);
nand g190(n898, n893, n799);
nand g191(n835, add2_i[28], n982);
nand g192(n856, n853, n858);
nand g193(n853, add1_i[25], n975);
or g194(n854, n975, add1_i[25]);
nand g195(n872, xenc27, n873);
nand g196(n878, add1_i[20], n881);
nand g197(n892, add2_i[17], n893);
nand g198(n926, n928, n929);
nand g199(n935, n933, xenc1);
nand g200(n809, n933, n801, xenc1);
nand g201(n811, n815, n936);
nand g202(result_o[32], xenc24, n822);
nand g203(n808, n994, n810);
nand g204(n860, add1_i[24], n863);
nand g205(n881, n883, n882);
nand g206(n883, add2_i[19], xenc56);
nand g207(n901, add1_i[16], n904);
nand g208(n904, n905, n906);
nand g209(n923, add1_i[11], n926);
nand g210(n932, add2_i[9], xenc12);
nand g211(n936, add2_i[7], n814);
nand g212(n955, add1_i[3], xenc10);
nand g213(n961, add1_i[1], n886);
or g214(n963, n886, add1_i[1]);
nand g215(n822, add2_i[31], n823);
nor g216(n895, xenc39, n897);
nand g217(n825, add1_i[30], xenc14);
not g218(n796, n991);
nand g219(n858, n859, add2_i[25]);
nand g220(n866, add2_i[23], n867);
nand g221(n870, add2_i[22], n871);
nand g222(n874, add2_i[21], n875);
nand g223(n882, xenc33, add1_i[19]);
not g224(n799, n897);
nand g225(n906, add2_i[15], n907);
nand g226(n909, add1_i[14], n912);
nand g227(n920, add2_i[12], xenc41);
nand g228(n929, add2_i[10], xenc53);
nand g229(n944, n984, n803, xenc9);
nand g230(n814, n984, n803, xenc11);
nand g231(n942, add1_i[7], n816, add2_i[6]);
or g232(n941, n984, n803);
nand g233(n953, n818, add2_i[4]);
nand g234(n959, add2_i[2], n837);
xor g235(xenc0, n862, keyinput0);
xor g236(xenc1, n934, keyinput1);
xor g237(result_o[1], xenc2, keyinput2);
xnor g238(xenc3, n878, keyinput3);
xor g239(xenc4, n870, keyinput4);
xnor g240(xenc5, n974, keyinput5);
xnor g241(xenc6, n962, keyinput6);
xor g242(xenc7, n942, keyinput7);
xnor g243(result_o[25], xenc8, keyinput8);
xor g244(xenc9, n945, keyinput9);
xor g245(xenc10, n819, keyinput10);
xor g246(xenc11, n938, keyinput11);
xnor g247(xenc12, n809, keyinput12);
xnor g248(xenc13, n845, keyinput13);
xor g249(xenc14, n828, keyinput14);
xor g250(xenc15, n946, keyinput15);
xor g251(xenc16, n972, keyinput16);
xnor g252(xenc17, n919, keyinput17);
xnor g253(xenc18, n856, keyinput18);
xor g254(xenc19, n895, keyinput19);
xnor g255(xenc20, n891, keyinput20);
xnor g256(xenc21, n922, keyinput21);
xnor g257(result_o[12], xenc22, keyinput22);
xor g258(result_o[22], xenc23, keyinput23);
xnor g259(xenc24, n821, keyinput24);
xnor g260(xenc25, n987, keyinput25);
xnor g261(result_o[21], xenc26, keyinput26);
xor g262(xenc27, n874, keyinput27);
xnor g263(xenc28, n965, keyinput28);
xor g264(xenc29, n854, keyinput29);
xnor g265(xenc30, n909, keyinput30);
xor g266(xenc31, n840, keyinput31);
xnor g267(xenc32, n887, keyinput32);
xor g268(xenc33, n885, keyinput33);
xor g269(xenc34, n868, keyinput34);
xor g270(xenc35, n927, keyinput35);
xnor g271(xenc36, n841, keyinput36);
xor g272(xenc37, n989, keyinput37);
xnor g273(result_o[26], xenc38, keyinput38);
xnor g274(xenc39, n896, keyinput39);
xnor g275(result_o[31], xenc40, keyinput40);
xor g276(xenc41, n921, keyinput41);
xor g277(xenc42, n820, keyinput42);
xor g278(xenc43, n957, keyinput43);
xor g279(xenc44, n797, keyinput44);
xnor g280(result_o[30], xenc45, keyinput45);
xnor g281(xenc46, n861, keyinput46);
xnor g282(xenc47, n808, keyinput47);
xor g283(result_o[2], xenc48, keyinput48);
xnor g284(xenc49, n824, keyinput49);
xor g285(xenc50, n920, keyinput50);
xor g286(xenc51, n943, keyinput51);
xnor g287(result_o[9], xenc52, keyinput52);
xnor g288(xenc53, n930, keyinput53);
xnor g289(result_o[20], xenc54, keyinput54);
xor g290(xenc55, n890, keyinput55);
xnor g291(xenc56, n884, keyinput56);
xnor g292(result_o[3], xenc57, keyinput57);
xnor g293(xenc58, n981, keyinput58);
xor g294(result_o[19], xenc59, keyinput59);
xor g295(xenc60, n961, keyinput60);
xnor g296(xenc61, n850, keyinput61);
xnor g297(xenc62, n1008, keyinput62);
xor g298(result_o[23], xenc63, keyinput63);
endmodule
