module carry_lookahead_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n655, n656, n658, n659, n660, n662, n663, n664, n665, n666, n668,
         n669, n670, n671, n672, n673, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n697, n698, n699, n700, n701, n702, n703, n705,
         n707, n708, n711, n712, n714, n715, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n739, n740, n742, n743, n744, n745,
         n747, n749, n750, n752, n753, n754, n755, n757, n759, n760, n761,
         n762, n763, n764, n765, n767, n769, n770, n772, n773, n774, n775,
         n777, n779, n780, n782, n783, n784, n785, n787, n788, n790, n791,
         n792, n793, n794, n795, n798, n799, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891;

  xor U672 ( result_o[8], n659, n660);
  xor U673 ( n660, add2_i[8], add1_i[8]);
  xor U674 ( result_o[6], n663, n664);
  xor U675 ( n664, add2_i[6], add1_i[6]);
  xor U676 ( result_o[5], n665, n666);
  xor U677 ( n666, add2_i[5], add1_i[5]);
  xor U678 ( result_o[3], n668, n669);
  xor U679 ( n669, add2_i[3], add1_i[3]);
  xor U680 ( result_o[30], n678, n679);
  xor U681 ( n679, add2_i[30], add1_i[30]);
  xor U682 ( result_o[2], n684, n685);
  xor U683 ( n685, add2_i[2], add1_i[2]);
  xor U684 ( result_o[28], n690, n691);
  xor U685 ( n691, add2_i[28], add1_i[28]);
  xor U686 ( result_o[26], n700, n701);
  xor U687 ( n701, add2_i[26], add1_i[26]);
  xor U688 ( result_o[24], n872, n711);
  xor U689 ( n711, add2_i[24], add1_i[24]);
  xor U690 ( result_o[22], n720, n721);
  xor U691 ( n721, add2_i[22], add1_i[22]);
  xor U692 ( result_o[20], n730, n731);
  xor U693 ( n731, add2_i[20], add1_i[20]);
  xor U694 ( result_o[1], n736, n737);
  xor U695 ( n737, add2_i[1], add1_i[1]);
  xor U696 ( result_o[18], n742, n743);
  xor U697 ( n743, add2_i[18], add1_i[18]);
  xor U698 ( result_o[16], n752, n753);
  xor U699 ( n753, add2_i[16], add1_i[16]);
  xor U700 ( result_o[14], n762, n763);
  xor U701 ( n763, add2_i[14], add1_i[14]);
  xor U702 ( result_o[12], n772, n773);
  xor U703 ( n773, add2_i[12], add1_i[12]);
  xor U704 ( result_o[10], n782, n783);
  xor U705 ( n783, add2_i[10], add1_i[10]);
  or U706 ( n736, add2_i[0], add1_i[0]);
  not U707 ( n830, add2_i[8]);
  not U708 ( n826, add2_i[12]);
  not U709 ( n832, add2_i[16]);
  not U710 ( n828, add2_i[9]);
  not U711 ( n836, add2_i[11]);
  not U712 ( n838, add2_i[17]);
  not U713 ( n834, add2_i[18]);
  nand U714 ( n665, n814, n815);
  nand U715 ( n814, add1_i[4], n803);
  nand U716 ( n815, add2_i[4], n802);
  or U717 ( n816, add2_i[0], add1_i[1]);
  or U718 ( n817, n827, n826);
  and U719 ( n889, n817, n818);
  and U720 ( n818, n819, n769);
  not U721 ( n819, add1_i[13]);
  or U722 ( n820, n833, n832);
  and U723 ( n839, n820, n821);
  and U724 ( n821, n822, n749);
  not U725 ( n822, add1_i[17]);
  or U726 ( n823, n831, n830);
  and U727 ( n829, n823, n824);
  and U728 ( n824, n825, n787);
  not U729 ( n825, add1_i[9]);
  or U730 ( n770, n826, n827);
  nor U731 ( n827, n772, add1_i[12]);
  or U732 ( n785, n829, n828);
  not U733 ( n864, add2_i[10]);
  or U734 ( n788, n830, n831);
  nor U735 ( n831, n659, add1_i[8]);
  or U736 ( n750, n832, n833);
  nor U737 ( n833, n752, add1_i[16]);
  or U738 ( n740, n834, n835);
  nor U739 ( n835, n742, add1_i[18]);
  not U740 ( n888, add2_i[13]);
  not U741 ( n890, add2_i[15]);
  not U742 ( n875, add2_i[25]);
  or U743 ( n775, n836, n837);
  nor U744 ( n837, n777, add1_i[11]);
  or U745 ( n745, n838, n839);
  xor U746 ( result_o[31], n840, n673);
  xor U747 ( n840, add1_i[31], add2_i[31]);
  xor U748 ( result_o[27], n841, n695);
  xor U749 ( n841, add1_i[27], add2_i[27]);
  xor U750 ( result_o[29], n842, n683);
  xor U751 ( n842, add1_i[29], add2_i[29]);
  xor U752 ( result_o[23], n843, n715);
  xor U753 ( n843, add1_i[23], add2_i[23]);
  xor U754 ( result_o[25], n844, n705);
  xor U755 ( n844, add1_i[25], add2_i[25]);
  not U756 ( n655, add1_i[4]);
  nor U757 ( n845, n846, n847);
  and U758 ( n846, add1_i[5], n802, add2_i[4]);
  and U759 ( n847, add1_i[5], n803, add1_i[4]);
  or U760 ( n729, n730, add1_i[20]);
  or U761 ( n799, n665, add1_i[5]);
  nor U762 ( n876, n848, n849);
  and U763 ( n848, n871, add2_i[24]);
  nand U764 ( n849, n861, n707);
  nor U765 ( n891, n850, n851);
  and U766 ( n850, n761, add2_i[14]);
  nand U767 ( n851, n860, n759);
  xor U768 ( result_o[17], n852, n747);
  xor U769 ( n852, add1_i[17], add2_i[17]);
  xor U770 ( result_o[19], n853, n735);
  xor U771 ( n853, add1_i[19], add2_i[19]);
  xor U772 ( result_o[15], n854, n757);
  xor U773 ( n854, add1_i[15], add2_i[15]);
  xnor U774 ( n726, add1_i[21], add2_i[21]);
  xor U775 ( result_o[13], n855, n767);
  xor U776 ( n855, add1_i[13], add2_i[13]);
  xor U777 ( result_o[9], n856, n658);
  xor U778 ( n856, add1_i[9], add2_i[9]);
  xor U779 ( result_o[11], n857, n777);
  xor U780 ( n857, add1_i[11], add2_i[11]);
  xor U781 ( result_o[7], n858, n662);
  xor U782 ( n858, add1_i[7], add2_i[7]);
  xor U783 ( result_o[4], n656, n859);
  xor U784 ( n859, add2_i[4], n655);
  not U785 ( n860, add1_i[15]);
  not U786 ( n861, add1_i[25]);
  nand U787 ( n714, n717, n862);
  and U788 ( n862, n718, n863);
  not U789 ( n863, add1_i[23]);
  or U790 ( n780, n865, n864);
  nor U791 ( n865, n782, add1_i[10]);
  nand U792 ( n866, n714, n869);
  and U793 ( n707, n866, n867);
  or U794 ( n867, n868, n712);
  not U795 ( n868, add1_i[24]);
  and U796 ( n869, add2_i[23], add1_i[24]);
  nand U797 ( n870, add2_i[23], n714);
  nand U798 ( n708, n871, add2_i[24]);
  nand U799 ( n871, n873, n874);
  nand U800 ( n872, n712, n870);
  nand U801 ( n873, n714, add2_i[23]);
  and U802 ( n874, n868, n712);
  or U803 ( n703, n876, n875);
  nand U804 ( n877, n729, n880);
  and U805 ( n722, n877, n878);
  or U806 ( n878, n879, n727);
  not U807 ( n879, add1_i[21]);
  and U808 ( n880, add2_i[20], add1_i[21]);
  nand U809 ( n881, n729, add2_i[20]);
  nand U810 ( n724, n881, n882);
  and U811 ( n882, n879, n727);
  nand U812 ( n725, n727, n728);
  nand U813 ( n805, add2_i[3], n806);
  nand U814 ( n792, n883, n793);
  and U815 ( n883, n794, n884);
  not U816 ( n884, add1_i[7]);
  nand U817 ( n662, n793, n794);
  nand U818 ( n885, n799, add2_i[5]);
  nand U819 ( n795, n885, n886);
  and U820 ( n886, n887, n845);
  not U821 ( n887, add1_i[6]);
  nand U822 ( n813, add2_i[0], add1_i[0]);
  nand U823 ( n663, n798, n845);
  nand U824 ( n676, add2_i[30], n677);
  nand U825 ( n798, n799, add2_i[5]);
  nand U826 ( n688, add2_i[28], n689);
  nand U827 ( n683, n687, n688);
  nand U828 ( n747, n749, n750);
  nand U829 ( n767, n769, n770);
  or U830 ( n765, n888, n889);
  or U831 ( n755, n890, n891);
  nand U832 ( n811, add2_i[1], n812);
  nand U833 ( n684, n810, n811);
  nand U834 ( n658, n787, n788);
  nand U835 ( n705, n707, n708);
  nand U836 ( result_o[32], n670, n671);
  nand U837 ( n695, n697, n698);
  nand U838 ( n718, add2_i[22], n719);
  nand U839 ( n727, add1_i[20], n730);
  nand U840 ( n760, add2_i[14], n761);
  nand U841 ( n769, add1_i[12], n772);
  nand U842 ( n787, add1_i[8], n659);
  nand U843 ( n794, add2_i[6], n795);
  nand U844 ( n804, add1_i[3], n668);
  or U845 ( n806, n668, add1_i[3]);
  nand U846 ( n807, add1_i[2], n684);
  or U847 ( n809, n684, add1_i[2]);
  nand U848 ( n728, add2_i[20], n729);
  nand U849 ( n671, add2_i[31], n672);
  nand U850 ( n698, add2_i[26], n699);
  nand U851 ( n700, n703, n702);
  nand U852 ( n752, n755, n754);
  nand U853 ( n668, n807, n808);
  nand U854 ( n808, add2_i[2], n809);
  nand U855 ( n730, n732, n733);
  nand U856 ( n733, add2_i[19], n734);
  nand U857 ( n772, n774, n775);
  nand U858 ( n659, n790, n791);
  nand U859 ( n791, n792, add2_i[7]);
  nand U860 ( n675, add1_i[30], n678);
  or U861 ( n677, n678, add1_i[30]);
  nand U862 ( n687, add1_i[28], n690);
  or U863 ( n689, n690, add1_i[28]);
  nand U864 ( n717, add1_i[22], n720);
  or U865 ( n719, n720, add1_i[22]);
  nand U866 ( n739, add1_i[18], n742);
  nand U867 ( n759, add1_i[14], n762);
  or U868 ( n761, n762, add1_i[14]);
  nand U869 ( n779, add1_i[10], n782);
  nand U870 ( n673, n675, n676);
  nand U871 ( n715, n717, n718);
  nand U872 ( n735, n739, n740);
  nand U873 ( n757, n759, n760);
  nand U874 ( n777, n780, n779);
  nand U875 ( n802, n656, n655);
  nand U876 ( n678, n680, n681);
  nand U877 ( n681, add2_i[29], n682);
  nand U878 ( n690, n692, n693);
  nand U879 ( n693, add2_i[27], n694);
  nand U880 ( n720, n722, n723);
  nand U881 ( n723, n724, add2_i[21]);
  nand U882 ( n742, n744, n745);
  nand U883 ( n762, n764, n765);
  nand U884 ( n782, n784, n785);
  nand U885 ( n803, n805, n804);
  nand U886 ( result_o[0], n736, n813);
  xnor U887 ( result_o[21], n726, n725);
  nand U888 ( n670, add1_i[31], n673);
  or U889 ( n672, n673, add1_i[31]);
  nand U890 ( n680, add1_i[29], n683);
  or U891 ( n682, n683, add1_i[29]);
  nand U892 ( n692, add1_i[27], n695);
  or U893 ( n694, n695, add1_i[27]);
  nand U894 ( n697, add1_i[26], n700);
  or U895 ( n699, n700, add1_i[26]);
  nand U896 ( n702, add1_i[25], n705);
  nand U897 ( n712, add1_i[23], n715);
  nand U898 ( n732, add1_i[19], n735);
  or U899 ( n734, n735, add1_i[19]);
  nand U900 ( n744, add1_i[17], n747);
  nand U901 ( n749, add1_i[16], n752);
  nand U902 ( n754, add1_i[15], n757);
  nand U903 ( n764, add1_i[13], n767);
  nand U904 ( n774, add1_i[11], n777);
  nand U905 ( n784, add1_i[9], n658);
  nand U906 ( n790, add1_i[7], n662);
  nand U907 ( n793, add1_i[6], n663);
  not U908 ( n656, n803);
  nand U909 ( n810, add1_i[1], n736);
  or U910 ( n812, n816, add1_i[0]);
endmodule
