// Verilog File 
module carry_lookahead_adder32_aor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n659, xenc8, n660, xenc127, n664, xenc34, xenc101, xenc96, n666, 
n668, n669, xenc104, n678, xenc126, xenc52, n679, xenc94, xenc123, xenc121, 
n685, n690, xenc62, xenc88, n691, xenc59, n701, xenc85, xenc115, n711, 
xenc7, n721, n730, xenc27, xenc54, n731, xenc116, n737, n742, n743, 
xenc4, xenc65, xenc107, xenc43, n753, n762, n763, xenc67, xenc12, xenc42, 
n773, n782, xenc29, n783, n736, n830, n826, n832, n828, n836, 
n838, n834, n814, n815, n665, n803, n802, n816, xenc11, xenc57, 
n817, xenc44, n889, n819, n769, n818, n833, xenc32, n820, xenc16, 
xenc10, n839, n822, n749, n821, xenc102, n823, xenc117, n829, xenc5, 
xenc47, n824, n825, n770, n827, xenc73, n785, n864, n788, n831, 
n750, xenc41, n835, n740, n888, n890, n875, xenc31, n837, n775, 
xenc77, xenc58, xenc120, n745, n840, n673, n841, xenc93, n842, n683, 
xenc19, n715, xenc113, n843, n844, n705, n655, n846, xenc72, n845, 
n847, n729, n799, xenc49, xenc66, n876, xenc60, n848, xenc106, n707, 
n849, n850, xenc84, n891, n761, n860, xenc15, n851, xenc28, n747, 
n852, xenc46, xenc20, n853, xenc33, n757, n854, n726, n855, n767, 
xenc108, xenc70, n658, n856, xenc99, xenc118, n857, xenc35, xenc81, xenc82, 
n858, xenc55, xenc45, xenc0, n859, n861, n717, xenc24, n714, xenc92, 
n863, n862, n865, n780, n869, n866, xenc18, xenc119, n868, n712, 
n867, n870, n708, xenc21, xenc112, n871, n872, n873, n874, xenc69, 
xenc39, n703, xenc51, n877, n878, n722, xenc48, n727, n879, n880, 
n881, xenc100, xenc124, n724, n882, xenc78, n725, xenc125, n805, n883, 
xenc122, n792, xenc37, xenc63, n884, n662, n885, xenc68, n795, xenc103, 
xenc23, n886, n887, n813, n798, n663, n677, n676, n689, n688, 
n687, xenc2, xenc110, n765, n755, xenc89, n811, xenc61, xenc83, n684, 
n670, n671, xenc75, xenc95, xenc26, n695, n719, n718, n760, n787, 
xenc114, n794, n804, n806, n807, n809, n728, xenc87, xenc98, n698, 
n702, n700, xenc40, xenc80, n752, xenc56, xenc86, xenc13, n808, xenc111, 
n733, n734, xenc25, xenc97, n772, xenc17, xenc91, xenc14, n791, n675, 
n739, n759, n779, xenc105, xenc76, n735, xenc3, xenc6, n777, xenc22, 
n681, xenc30, xenc36, n693, xenc53, xenc9, xenc74, n720, n723, xenc50, 
xenc109, n764, xenc64, xenc38, xenc1, xenc90, xenc79, xenc71, n672, n680, 
n682, n692, n694, n697, n699, n732, n744, n754, n774, n784, 
n790, n793, n656, n810, n812;

xor g0(result_o[8], n659, xenc8);
xor g1(n660, add2_i[8], add1_i[8]);
xor g2(xenc34, xenc127, n664);
xor g3(n664, add2_i[6], add1_i[6]);
xor g4(result_o[5], xenc101, xenc96);
xor g5(n666, add2_i[5], add1_i[5]);
xor g6(xenc104, n668, n669);
xor g7(n669, add2_i[3], add1_i[3]);
xor g8(xenc52, n678, xenc126);
xor g9(n679, add2_i[30], add1_i[30]);
xor g10(xenc121, xenc94, xenc123);
xor g11(n685, add2_i[2], add1_i[2]);
xor g12(xenc88, n690, xenc62);
xor g13(n691, add2_i[28], add1_i[28]);
xor g14(xenc85, xenc59, n701);
xor g15(n701, add2_i[26], add1_i[26]);
xor g16(result_o[24], xenc115, n711);
xor g17(n711, add2_i[24], add1_i[24]);
xor g18(result_o[22], xenc7, n721);
xor g19(n721, add2_i[22], add1_i[22]);
xor g20(xenc54, n730, xenc27);
xor g21(n731, add2_i[20], add1_i[20]);
xor g22(result_o[1], xenc116, n737);
xor g23(n737, add2_i[1], add1_i[1]);
xor g24(xenc4, n742, n743);
xor g25(n743, add2_i[18], add1_i[18]);
xor g26(xenc43, xenc65, xenc107);
xor g27(n753, add2_i[16], add1_i[16]);
xor g28(result_o[14], n762, n763);
xor g29(n763, add2_i[14], add1_i[14]);
xor g30(xenc42, xenc67, xenc12);
xor g31(n773, add2_i[12], add1_i[12]);
xor g32(result_o[10], n782, xenc29);
xor g33(n783, add2_i[10], add1_i[10]);
or g34(n736, add2_i[0], add1_i[0]);
not g35(n830, add2_i[8]);
not g36(n826, add2_i[12]);
not g37(n832, add2_i[16]);
not g38(n828, add2_i[9]);
not g39(n836, add2_i[11]);
not g40(n838, add2_i[17]);
not g41(n834, add2_i[18]);
nand g42(n665, n814, n815);
nand g43(n814, add1_i[4], n803);
nand g44(n815, add2_i[4], n802);
or g45(n816, add2_i[0], add1_i[1]);
or g46(n817, xenc11, xenc57);
and g47(n889, n817, xenc44);
and g48(n818, n819, n769);
not g49(n819, add1_i[13]);
or g50(n820, n833, xenc32);
and g51(n839, xenc16, xenc10);
and g52(n821, n822, n749);
not g53(n822, add1_i[17]);
or g54(n823, xenc102, n830);
and g55(n829, n823, xenc117);
and g56(n824, xenc5, xenc47);
not g57(n825, add1_i[9]);
or g58(n770, xenc57, xenc11);
nor g59(n827, xenc67, add1_i[12]);
or g60(n785, n829, xenc73);
not g61(n864, add2_i[10]);
or g62(n788, n830, xenc102);
nor g63(n831, n659, add1_i[8]);
or g64(n750, xenc32, n833);
nor g65(n833, xenc65, add1_i[16]);
or g66(n740, xenc41, n835);
nor g67(n835, n742, add1_i[18]);
not g68(n888, add2_i[13]);
not g69(n890, add2_i[15]);
not g70(n875, add2_i[25]);
or g71(n775, xenc31, n837);
nor g72(n837, xenc77, add1_i[11]);
or g73(n745, xenc58, xenc120);
xor g74(result_o[31], n840, n673);
xor g75(n840, add1_i[31], add2_i[31]);
xor g76(result_o[27], n841, xenc93);
xor g77(n841, add1_i[27], add2_i[27]);
xor g78(result_o[29], n842, n683);
xor g79(n842, add1_i[29], add2_i[29]);
xor g80(xenc113, xenc19, n715);
xor g81(n843, add1_i[23], add2_i[23]);
xor g82(result_o[25], n844, n705);
xor g83(n844, add1_i[25], add2_i[25]);
not g84(n655, add1_i[4]);
nor g85(n845, n846, xenc72);
and g86(n846, add1_i[5], n802, add2_i[4]);
and g87(n847, add1_i[5], n803, add1_i[4]);
or g88(n729, n730, add1_i[20]);
or g89(n799, xenc101, add1_i[5]);
nor g90(n876, xenc49, xenc66);
and g91(n848, xenc60, add2_i[24]);
nand g92(n849, xenc106, n707);
nor g93(n891, n850, xenc84);
and g94(n850, n761, add2_i[14]);
nand g95(n851, n860, xenc15);
xor g96(result_o[17], xenc28, n747);
xor g97(n852, add1_i[17], add2_i[17]);
xor g98(result_o[19], xenc46, xenc20);
xor g99(n853, add1_i[19], add2_i[19]);
xor g100(result_o[15], xenc33, n757);
xor g101(n854, add1_i[15], add2_i[15]);
xnor g102(n726, add1_i[21], add2_i[21]);
xor g103(xenc108, n855, n767);
xor g104(n855, add1_i[13], add2_i[13]);
xor g105(result_o[9], xenc70, n658);
xor g106(n856, add1_i[9], add2_i[9]);
xor g107(xenc118, xenc99, xenc77);
xor g108(n857, add1_i[11], add2_i[11]);
xor g109(xenc82, xenc35, xenc81);
xor g110(n858, add1_i[7], add2_i[7]);
xor g111(xenc0, xenc55, xenc45);
xor g112(n859, add2_i[4], n655);
not g113(n860, add1_i[15]);
not g114(n861, add1_i[25]);
nand g115(n714, n717, xenc24);
and g116(n862, xenc92, n863);
not g117(n863, add1_i[23]);
or g118(n780, n865, n864);
nor g119(n865, n782, add1_i[10]);
nand g120(n866, n714, n869);
and g121(n707, xenc18, xenc119);
or g122(n867, n868, n712);
not g123(n868, add1_i[24]);
and g124(n869, add2_i[23], add1_i[24]);
nand g125(n870, add2_i[23], n714);
nand g126(n708, xenc60, add2_i[24]);
nand g127(n871, xenc21, xenc112);
nand g128(n872, n712, n870);
nand g129(n873, n714, add2_i[23]);
and g130(n874, n868, n712);
or g131(n703, xenc69, xenc39);
nand g132(n877, n729, xenc51);
and g133(n722, n877, n878);
or g134(n878, xenc48, n727);
not g135(n879, add1_i[21]);
and g136(n880, add2_i[20], add1_i[21]);
nand g137(n881, n729, add2_i[20]);
nand g138(n724, xenc100, xenc124);
and g139(n882, xenc48, n727);
nand g140(n725, n727, xenc78);
nand g141(n805, add2_i[3], xenc125);
nand g142(n792, n883, xenc122);
and g143(n883, xenc37, xenc63);
not g144(n884, add1_i[7]);
nand g145(n662, xenc122, xenc37);
nand g146(n885, n799, add2_i[5]);
nand g147(n795, n885, xenc68);
and g148(n886, xenc103, xenc23);
not g149(n887, add1_i[6]);
nand g150(n813, add2_i[0], add1_i[0]);
nand g151(n663, n798, xenc23);
nand g152(n676, add2_i[30], n677);
nand g153(n798, n799, add2_i[5]);
nand g154(n688, add2_i[28], n689);
nand g155(n683, n687, xenc2);
nand g156(n747, n749, n750);
nand g157(n767, n769, n770);
or g158(n765, n888, xenc110);
or g159(n755, n890, n891);
nand g160(n811, add2_i[1], xenc89);
nand g161(n684, xenc61, xenc83);
nand g162(n658, xenc47, n788);
nand g163(n705, n707, n708);
nand g164(xenc75, n670, n671);
nand g165(n695, xenc95, xenc26);
nand g166(n718, add2_i[22], n719);
nand g167(n727, add1_i[20], n730);
nand g168(n760, add2_i[14], n761);
nand g169(n769, add1_i[12], xenc67);
nand g170(n787, add1_i[8], n659);
nand g171(n794, add2_i[6], xenc114);
nand g172(n804, add1_i[3], n668);
or g173(n806, n668, add1_i[3]);
nand g174(n807, add1_i[2], xenc94);
or g175(n809, xenc94, add1_i[2]);
nand g176(n728, add2_i[20], n729);
nand g177(n671, add2_i[31], xenc87);
nand g178(n698, add2_i[26], xenc98);
nand g179(n700, n703, n702);
nand g180(n752, xenc40, xenc80);
nand g181(n668, xenc56, xenc86);
nand g182(n808, add2_i[2], xenc13);
nand g183(n730, xenc111, n733);
nand g184(n733, add2_i[19], n734);
nand g185(n772, xenc25, xenc97);
nand g186(n659, xenc17, xenc91);
nand g187(n791, xenc14, add2_i[7]);
nand g188(n675, add1_i[30], n678);
or g189(n677, n678, add1_i[30]);
nand g190(n687, add1_i[28], n690);
or g191(n689, n690, add1_i[28]);
nand g192(n717, add1_i[22], xenc7);
or g193(n719, xenc7, add1_i[22]);
nand g194(n739, add1_i[18], n742);
nand g195(n759, add1_i[14], n762);
or g196(n761, n762, add1_i[14]);
nand g197(n779, add1_i[10], n782);
nand g198(n673, xenc105, n676);
nand g199(n715, n717, xenc92);
nand g200(n735, n739, xenc76);
nand g201(n757, xenc15, n760);
nand g202(n777, xenc3, xenc6);
nand g203(n802, xenc55, n655);
nand g204(n678, xenc22, n681);
nand g205(n681, add2_i[29], xenc30);
nand g206(n690, xenc36, n693);
nand g207(n693, add2_i[27], xenc53);
nand g208(n720, xenc9, xenc74);
nand g209(n723, n724, add2_i[21]);
nand g210(n742, xenc50, xenc109);
nand g211(n762, n764, xenc64);
nand g212(n782, xenc38, n785);
nand g213(n803, xenc1, n804);
nand g214(xenc90, xenc116, n813);
xnor g215(xenc71, n726, xenc79);
nand g216(n670, add1_i[31], n673);
or g217(n672, n673, add1_i[31]);
nand g218(n680, add1_i[29], n683);
or g219(n682, n683, add1_i[29]);
nand g220(n692, add1_i[27], xenc93);
or g221(n694, xenc93, add1_i[27]);
nand g222(n697, add1_i[26], xenc59);
or g223(n699, xenc59, add1_i[26]);
nand g224(n702, add1_i[25], n705);
nand g225(n712, add1_i[23], n715);
nand g226(n732, add1_i[19], xenc20);
or g227(n734, xenc20, add1_i[19]);
nand g228(n744, add1_i[17], n747);
nand g229(n749, add1_i[16], xenc65);
nand g230(n754, add1_i[15], n757);
nand g231(n764, add1_i[13], n767);
nand g232(n774, add1_i[11], xenc77);
nand g233(n784, add1_i[9], n658);
nand g234(n790, add1_i[7], xenc81);
nand g235(n793, add1_i[6], xenc127);
not g236(n656, n803);
nand g237(n810, add1_i[1], xenc116);
or g238(n812, n816, add1_i[0]);
or g239(result_o[4], xenc0, keyinput0);
or g240(xenc1, n805, keyinput1);
and g241(xenc2, n688, keyinput2);
or g242(xenc3, n780, keyinput3);
and g243(result_o[18], xenc4, keyinput4);
or g244(xenc5, n825, keyinput5);
or g245(xenc6, n779, keyinput6);
and g246(xenc7, n720, keyinput7);
or g247(xenc8, n660, keyinput8);
and g248(xenc9, n722, keyinput9);
or g249(xenc10, n821, keyinput10);
and g250(xenc11, n827, keyinput11);
and g251(xenc12, n773, keyinput12);
and g252(xenc13, n809, keyinput13);
or g253(xenc14, n792, keyinput14);
or g254(xenc15, n759, keyinput15);
and g255(xenc16, n820, keyinput16);
or g256(xenc17, n790, keyinput17);
and g257(xenc18, n866, keyinput18);
and g258(xenc19, n843, keyinput19);
and g259(xenc20, n735, keyinput20);
or g260(xenc21, n873, keyinput21);
or g261(xenc22, n680, keyinput22);
and g262(xenc23, n845, keyinput23);
or g263(xenc24, n862, keyinput24);
or g264(xenc25, n774, keyinput25);
and g265(xenc26, n698, keyinput26);
or g266(xenc27, n731, keyinput27);
and g267(xenc28, n852, keyinput28);
or g268(xenc29, n783, keyinput29);
and g269(xenc30, n682, keyinput30);
or g270(xenc31, n836, keyinput31);
and g271(xenc32, n832, keyinput32);
and g272(xenc33, n854, keyinput33);
or g273(result_o[6], xenc34, keyinput34);
and g274(xenc35, n858, keyinput35);
and g275(xenc36, n692, keyinput36);
and g276(xenc37, n794, keyinput37);
and g277(xenc38, n784, keyinput38);
or g278(xenc39, n875, keyinput39);
and g279(xenc40, n755, keyinput40);
or g280(xenc41, n834, keyinput41);
or g281(result_o[12], xenc42, keyinput42);
and g282(result_o[16], xenc43, keyinput43);
or g283(xenc44, n818, keyinput44);
and g284(xenc45, n859, keyinput45);
and g285(xenc46, n853, keyinput46);
or g286(xenc47, n787, keyinput47);
or g287(xenc48, n879, keyinput48);
and g288(xenc49, n848, keyinput49);
and g289(xenc50, n744, keyinput50);
or g290(xenc51, n880, keyinput51);
or g291(result_o[30], xenc52, keyinput52);
or g292(xenc53, n694, keyinput53);
and g293(result_o[20], xenc54, keyinput54);
and g294(xenc55, n656, keyinput55);
or g295(xenc56, n807, keyinput56);
and g296(xenc57, n826, keyinput57);
and g297(xenc58, n838, keyinput58);
or g298(xenc59, n700, keyinput59);
or g299(xenc60, n871, keyinput60);
and g300(xenc61, n810, keyinput61);
or g301(xenc62, n691, keyinput62);
or g302(xenc63, n884, keyinput63);
and g303(xenc64, n765, keyinput64);
and g304(xenc65, n752, keyinput65);
or g305(xenc66, n849, keyinput66);
and g306(xenc67, n772, keyinput67);
and g307(xenc68, n886, keyinput68);
or g308(xenc69, n876, keyinput69);
or g309(xenc70, n856, keyinput70);
and g310(result_o[21], xenc71, keyinput71);
and g311(xenc72, n847, keyinput72);
and g312(xenc73, n828, keyinput73);
and g313(xenc74, n723, keyinput74);
or g314(result_o[32], xenc75, keyinput75);
and g315(xenc76, n740, keyinput76);
and g316(xenc77, n777, keyinput77);
and g317(xenc78, n728, keyinput78);
or g318(xenc79, n725, keyinput79);
and g319(xenc80, n754, keyinput80);
and g320(xenc81, n662, keyinput81);
or g321(result_o[7], xenc82, keyinput82);
and g322(xenc83, n811, keyinput83);
and g323(xenc84, n851, keyinput84);
or g324(result_o[26], xenc85, keyinput85);
and g325(xenc86, n808, keyinput86);
or g326(xenc87, n672, keyinput87);
or g327(result_o[28], xenc88, keyinput88);
and g328(xenc89, n812, keyinput89);
and g329(result_o[0], xenc90, keyinput90);
and g330(xenc91, n791, keyinput91);
and g331(xenc92, n718, keyinput92);
or g332(xenc93, n695, keyinput93);
or g333(xenc94, n684, keyinput94);
or g334(xenc95, n697, keyinput95);
or g335(xenc96, n666, keyinput96);
and g336(xenc97, n775, keyinput97);
or g337(xenc98, n699, keyinput98);
or g338(xenc99, n857, keyinput99);
or g339(xenc100, n881, keyinput100);
or g340(xenc101, n665, keyinput101);
or g341(xenc102, n831, keyinput102);
or g342(xenc103, n887, keyinput103);
or g343(result_o[3], xenc104, keyinput104);
and g344(xenc105, n675, keyinput105);
and g345(xenc106, n861, keyinput106);
and g346(xenc107, n753, keyinput107);
and g347(result_o[13], xenc108, keyinput108);
and g348(xenc109, n745, keyinput109);
or g349(xenc110, n889, keyinput110);
or g350(xenc111, n732, keyinput111);
or g351(xenc112, n874, keyinput112);
and g352(result_o[23], xenc113, keyinput113);
or g353(xenc114, n795, keyinput114);
or g354(xenc115, n872, keyinput115);
or g355(xenc116, n736, keyinput116);
or g356(xenc117, n824, keyinput117);
and g357(result_o[11], xenc118, keyinput118);
and g358(xenc119, n867, keyinput119);
and g359(xenc120, n839, keyinput120);
and g360(result_o[2], xenc121, keyinput121);
and g361(xenc122, n793, keyinput122);
and g362(xenc123, n685, keyinput123);
and g363(xenc124, n882, keyinput124);
or g364(xenc125, n806, keyinput125);
or g365(xenc126, n679, keyinput126);
or g366(xenc127, n663, keyinput127);
endmodule
