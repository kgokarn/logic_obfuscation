// Verilog File 
module error_tolerant_type2_adder32_aor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire xenc15, xenc39, n145, xenc65, xenc67, n146, n149, xenc16, n153, 
xenc8, n154, xenc40, xenc33, xenc10, n157, n171, xenc45, xenc80, n172, 
n188, xenc14, n189, n192, xenc49, n193, n175, xenc88, n176, xenc35, 
xenc119, xenc37, n196, n204, xenc44, n205, n217, xenc7, xenc6, n218, 
xenc9, n222, n221, xenc56, xenc114, xenc93, n225, n229, xenc122, xenc22, 
xenc92, n243, xenc85, xenc127, xenc53, n246, xenc124, xenc111, xenc82, n250, 
xenc107, xenc86, n255, n254, xenc36, n200, n201, xenc71, xenc47, n268, 
n271, xenc77, xenc99, xenc75, n276, n275, xenc5, xenc55, n279, xenc81, 
n293, xenc60, xenc2, n297, n296, n300, xenc42, n301, n304, xenc11, 
xenc57, xenc109, xenc27, n318, n321, xenc103, n322, n325, n143, n328, 
n144, n170, n142, xenc121, xenc115, n317, n319, n148, n295, n270, 
n245, n220, n191, n320, n155, xenc17, n156, xenc108, n303, n302, 
n277, n278, n252, n253, n251, xenc54, xenc90, n226, n227, n228, 
n202, n203, n197, n151, xenc51, n150, n152, xenc64, n299, n298, 
n273, xenc41, n272, n274, xenc94, xenc26, n247, n248, n249, n223, 
xenc91, n224, n194, xenc78, n195, xenc19, xenc83, n326, n327, n323, 
n324, xenc117, xenc70, xenc50, n329, n331, n330, n306, xenc74, n305, 
xenc13, n308, n307, xenc101, n282, n280, xenc0, n281, n283, xenc126, 
xenc72, xenc87, n256, xenc32, n257, n258, n231, xenc58, n230, xenc105, 
xenc18, n232, n233, xenc61, xenc34, n209, n206, n208, n207, n337, 
xenc123, n336, n339, n338, n314, xenc24, n313, xenc97, n315, n316, 
n289, n290, n288, n291, n264, n265, n263, n266, xenc100, xenc12, 
n238, n239, xenc59, n240, n241, xenc89, n215, n213, n214, xenc52, 
n216, xenc38, n164, n162, xenc112, n163, xenc63, n165, xenc76, n334, 
n332, xenc116, n333, xenc46, n335, xenc95, xenc25, n309, n310, xenc21, 
n311, n312, xenc43, xenc3, n284, xenc28, n285, xenc79, n286, n287, 
xenc125, xenc20, n259, n260, xenc106, n261, n262, n235, n236, n234, 
xenc4, xenc118, n237, n210, xenc69, xenc31, n212, n211, n159, n160, 
n158, n161, n147, n294, n292, xenc1, xenc23, n267, n269, n244, 
xenc30, n242, n219, xenc96, xenc68, n190, xenc104, n168, n166, xenc110, 
n167, xenc113, n169, n173, xenc62, n174, xenc84, xenc120, n199, n198, 
n185, n186, n184, n187, xenc98, n182, n180, xenc48, n181, xenc29, 
n183, xenc73, xenc102, xenc66, n177, n179, n178;

xor g0(result_o[9], xenc15, add2_i[9]);
xor g1(result_o[8], xenc39, add2_i[8]);
xor g2(xenc67, n145, xenc65);
xor g3(n146, add2_i[7], add1_i[7]);
xor g4(result_o[6], add2_i[6], n149);
xor g5(n149, xenc16, add1_i[6]);
xor g6(xenc8, n153, add2_i[5]);
xor g7(n153, n154, add1_i[5]);
xor g8(xenc33, xenc40, add2_i[4]);
xor g9(n157, xenc10, add1_i[4]);
xor g10(xenc80, n171, xenc45);
xor g11(n172, add2_i[3], add1_i[3]);
xor g12(result_o[31], n188, xenc14);
xor g13(n189, add2_i[31], add1_i[31]);
xor g14(xenc49, add2_i[30], n192);
xor g15(n192, n193, add1_i[30]);
xor g16(xenc88, add2_i[2], n175);
xor g17(n175, n176, add1_i[2]);
xor g18(xenc119, xenc35, add2_i[29]);
xor g19(n196, xenc37, add1_i[29]);
xor g20(xenc44, n204, add2_i[28]);
xor g21(n204, n205, add1_i[28]);
xor g22(xenc6, n217, xenc7);
xor g23(n218, add2_i[27], add1_i[27]);
xor g24(result_o[26], add2_i[26], xenc9);
xor g25(n221, n222, add1_i[26]);
xor g26(xenc114, xenc56, add2_i[25]);
xor g27(n225, xenc93, add1_i[25]);
xor g28(xenc122, n229, add2_i[24]);
xor g29(n229, xenc22, add1_i[24]);
xor g30(xenc85, xenc92, n243);
xor g31(n243, add2_i[23], add1_i[23]);
xor g32(result_o[22], add2_i[22], xenc127);
xor g33(n246, xenc53, add1_i[22]);
xor g34(xenc111, xenc124, add2_i[21]);
xor g35(n250, xenc82, add1_i[21]);
xor g36(xenc86, xenc107, add2_i[20]);
xor g37(n254, n255, add1_i[20]);
xor g38(result_o[1], xenc36, add2_i[1]);
xor g39(n201, n200, add1_i[1]);
xor g40(result_o[19], xenc71, xenc47);
xor g41(n268, add2_i[19], add1_i[19]);
xor g42(xenc77, add2_i[18], n271);
xor g43(n271, xenc99, add1_i[18]);
xor g44(result_o[17], xenc75, add2_i[17]);
xor g45(n275, n276, add1_i[17]);
xor g46(result_o[16], xenc5, add2_i[16]);
xor g47(n279, xenc55, add1_i[16]);
xor g48(xenc60, xenc81, n293);
xor g49(n293, add2_i[15], add1_i[15]);
xor g50(result_o[14], add2_i[14], xenc2);
xor g51(n296, n297, add1_i[14]);
xor g52(xenc42, n300, add2_i[13]);
xor g53(n300, n301, add1_i[13]);
xor g54(result_o[12], n304, add2_i[12]);
xor g55(n304, xenc11, add1_i[12]);
xor g56(xenc27, xenc57, xenc109);
xor g57(n318, add2_i[11], add1_i[11]);
xor g58(xenc103, n321, add2_i[10]);
xor g59(n321, n322, add1_i[10]);
xor g60(n143, n325, add1_i[9]);
xor g61(n144, n328, add1_i[8]);
not g62(n142, n170);
nand g63(result_o[0], n170, n200);
nand g64(n317, xenc121, xenc115);
nand g65(n319, add1_i[10], n322);
nand g66(n148, n149, add2_i[6]);
nand g67(n295, xenc2, add2_i[14]);
nand g68(n270, n271, add2_i[18]);
nand g69(n245, xenc127, add2_i[22]);
nand g70(n220, xenc9, add2_i[26]);
nand g71(n191, n192, add2_i[30]);
nand g72(n320, n321, add2_i[10]);
nand g73(n170, add2_i[0], add1_i[0]);
nand g74(n154, n155, xenc17);
nand g75(n155, add1_i[4], xenc10);
nand g76(n156, xenc40, add2_i[4]);
nand g77(n301, xenc108, n303);
nand g78(n302, add1_i[12], xenc11);
nand g79(n303, n304, add2_i[12]);
nand g80(n276, n277, n278);
nand g81(n277, add1_i[16], xenc55);
nand g82(n278, xenc5, add2_i[16]);
nand g83(n251, n252, n253);
nand g84(n252, add1_i[20], n255);
nand g85(n253, xenc107, add2_i[20]);
nand g86(n226, xenc54, xenc90);
nand g87(n227, add1_i[24], xenc22);
nand g88(n228, n229, add2_i[24]);
nand g89(n197, n202, n203);
nand g90(n202, add1_i[28], n205);
nand g91(n203, n204, add2_i[28]);
nand g92(n150, n151, xenc51);
nand g93(n151, add1_i[5], n154);
nand g94(n152, n153, add2_i[5]);
nand g95(n297, xenc64, n299);
nand g96(n298, add1_i[13], n301);
nand g97(n299, n300, add2_i[13]);
nand g98(n272, n273, xenc41);
nand g99(n273, add1_i[17], n276);
nand g100(n274, xenc75, add2_i[17]);
nand g101(n247, xenc94, xenc26);
nand g102(n248, add1_i[21], xenc82);
nand g103(n249, xenc124, add2_i[21]);
nand g104(n222, n223, xenc91);
nand g105(n223, add1_i[25], xenc93);
nand g106(n224, xenc56, add2_i[25]);
nand g107(n193, n194, xenc78);
nand g108(n194, add1_i[29], xenc37);
nand g109(n195, xenc35, add2_i[29]);
nand g110(n325, xenc19, xenc83);
nand g111(n326, add1_i[8], n328);
nand g112(n327, add2_i[8], xenc39);
nand g113(n322, n323, n324);
nand g114(n323, add1_i[9], n325);
nand g115(n324, add2_i[9], xenc15);
nand g116(n328, xenc117, xenc70);
nand g117(n329, add1_i[7], xenc50);
nand g118(n330, add2_i[7], n331);
or g119(n331, xenc50, add1_i[7]);
nand g120(n305, n306, xenc74);
nand g121(n306, add1_i[11], xenc13);
nand g122(n307, add2_i[11], n308);
or g123(n308, xenc13, add1_i[11]);
nand g124(n280, xenc101, n282);
nand g125(n281, add1_i[15], xenc0);
nand g126(n282, add2_i[15], n283);
or g127(n283, xenc0, add1_i[15]);
nand g128(n255, xenc126, xenc72);
nand g129(n256, add1_i[19], xenc87);
nand g130(n257, add2_i[19], xenc32);
or g131(n258, xenc87, add1_i[19]);
nand g132(n230, n231, xenc58);
nand g133(n231, add1_i[23], xenc105);
nand g134(n232, add2_i[23], xenc18);
or g135(n233, xenc105, add1_i[23]);
nand g136(n205, xenc61, xenc34);
nand g137(n206, add1_i[27], n209);
nand g138(n207, add2_i[27], n208);
or g139(n208, n209, add1_i[27]);
nand g140(n336, n337, xenc123);
nand g141(n337, add2_i[5], add1_i[5]);
nand g142(n338, add1_i[4], n339, add2_i[4]);
or g143(n339, add2_i[5], add1_i[5]);
nand g144(n313, n314, xenc24);
nand g145(n314, add2_i[9], add1_i[9]);
nand g146(n315, add1_i[8], xenc97, add2_i[8]);
or g147(n316, add2_i[9], add1_i[9]);
nand g148(n288, n289, n290);
nand g149(n289, add2_i[13], add1_i[13]);
nand g150(n290, add1_i[12], n291, add2_i[12]);
or g151(n291, add2_i[13], add1_i[13]);
nand g152(n263, n264, n265);
nand g153(n264, add2_i[17], add1_i[17]);
nand g154(n265, add1_i[16], n266, add2_i[16]);
or g155(n266, add2_i[17], add1_i[17]);
nand g156(n238, xenc100, xenc12);
nand g157(n239, add2_i[21], add1_i[21]);
nand g158(n240, add1_i[20], xenc59, add2_i[20]);
or g159(n241, add2_i[21], add1_i[21]);
nand g160(n213, xenc89, n215);
nand g161(n214, add2_i[25], add1_i[25]);
nand g162(n215, add1_i[24], xenc52, add2_i[24]);
or g163(n216, add2_i[25], add1_i[25]);
nand g164(n162, xenc38, n164);
nand g165(n163, add1_i[2], xenc112);
nand g166(n164, add2_i[2], xenc63);
or g167(n165, xenc112, add1_i[2]);
nand g168(n332, xenc76, n334);
nand g169(n333, add1_i[6], xenc116);
nand g170(n334, add2_i[6], xenc46);
or g171(n335, xenc116, add1_i[6]);
nand g172(n309, xenc95, xenc25);
nand g173(n310, add1_i[10], n313);
nand g174(n311, add2_i[10], xenc21);
or g175(n312, n313, add1_i[10]);
nand g176(n284, xenc43, xenc3);
nand g177(n285, add1_i[14], xenc28);
nand g178(n286, add2_i[14], xenc79);
or g179(n287, xenc28, add1_i[14]);
nand g180(n259, xenc125, xenc20);
nand g181(n260, add1_i[18], n263);
nand g182(n261, add2_i[18], xenc106);
or g183(n262, n263, add1_i[18]);
nand g184(n234, n235, n236);
nand g185(n235, add1_i[22], xenc4);
nand g186(n236, add2_i[22], xenc118);
or g187(n237, xenc4, add1_i[22]);
nand g188(n209, n210, xenc69);
nand g189(n210, add1_i[26], xenc31);
nand g190(n211, add2_i[26], n212);
or g191(n212, xenc31, add1_i[26]);
nand g192(n158, n159, n160);
nand g193(n159, add1_i[3], n162);
nand g194(n160, add2_i[3], n161);
or g195(n161, n162, add1_i[3]);
nand g196(n145, n147, n148);
nand g197(n147, add1_i[6], xenc16);
nand g198(n292, n294, n295);
nand g199(n294, add1_i[14], n297);
nand g200(n267, xenc1, xenc23);
nand g201(n269, add1_i[18], xenc99);
nand g202(n242, n244, xenc30);
nand g203(n244, add1_i[22], xenc53);
nand g204(n217, n219, xenc96);
nand g205(n219, add1_i[26], n222);
nand g206(n188, xenc68, n191);
nand g207(n190, add1_i[30], n193);
nand g208(n166, xenc104, n168);
nand g209(n167, add1_i[1], xenc110);
nand g210(n168, add2_i[1], xenc113);
or g211(n169, add1_i[1], xenc110);
or g212(n200, add2_i[0], add1_i[0]);
nand g213(n171, n173, xenc62);
nand g214(n173, add1_i[2], n176);
nand g215(n174, n175, add2_i[2]);
nand g216(n176, xenc84, xenc120);
nand g217(n199, add1_i[1], n200);
nand g218(n198, xenc36, add2_i[1]);
nand g219(n184, n185, n186);
nand g220(n185, add2_i[29], add1_i[29]);
nand g221(n186, add1_i[28], n187, add2_i[28]);
or g222(n187, add2_i[29], add1_i[29]);
nand g223(n180, xenc98, n182);
nand g224(n181, add1_i[30], xenc48);
nand g225(n182, add2_i[30], xenc29);
or g226(n183, xenc48, add1_i[30]);
nand g227(result_o[32], xenc73, xenc102);
nand g228(n177, add1_i[31], xenc66);
nand g229(n178, add2_i[31], n179);
or g230(n179, xenc66, add1_i[31]);
and g231(xenc0, n284, keyinput0);
or g232(xenc1, n269, keyinput1);
or g233(xenc2, n296, keyinput2);
or g234(xenc3, n286, keyinput3);
or g235(xenc4, n238, keyinput4);
or g236(xenc5, n279, keyinput5);
or g237(result_o[27], xenc6, keyinput6);
and g238(xenc7, n218, keyinput7);
or g239(result_o[5], xenc8, keyinput8);
and g240(xenc9, n221, keyinput9);
and g241(xenc10, n158, keyinput10);
and g242(xenc11, n305, keyinput11);
or g243(xenc12, n240, keyinput12);
or g244(xenc13, n309, keyinput13);
and g245(xenc14, n189, keyinput14);
and g246(xenc15, n143, keyinput15);
or g247(xenc16, n150, keyinput16);
or g248(xenc17, n156, keyinput17);
or g249(xenc18, n233, keyinput18);
or g250(xenc19, n326, keyinput19);
and g251(xenc20, n261, keyinput20);
or g252(xenc21, n312, keyinput21);
and g253(xenc22, n230, keyinput22);
and g254(xenc23, n270, keyinput23);
or g255(xenc24, n315, keyinput24);
or g256(xenc25, n311, keyinput25);
and g257(xenc26, n249, keyinput26);
or g258(result_o[11], xenc27, keyinput27);
and g259(xenc28, n288, keyinput28);
and g260(xenc29, n183, keyinput29);
and g261(xenc30, n245, keyinput30);
and g262(xenc31, n213, keyinput31);
or g263(xenc32, n258, keyinput32);
or g264(result_o[4], xenc33, keyinput33);
or g265(xenc34, n207, keyinput34);
and g266(xenc35, n196, keyinput35);
and g267(xenc36, n201, keyinput36);
and g268(xenc37, n197, keyinput37);
or g269(xenc38, n163, keyinput38);
and g270(xenc39, n144, keyinput39);
and g271(xenc40, n157, keyinput40);
or g272(xenc41, n274, keyinput41);
and g273(result_o[13], xenc42, keyinput42);
or g274(xenc43, n285, keyinput43);
and g275(result_o[28], xenc44, keyinput44);
or g276(xenc45, n172, keyinput45);
or g277(xenc46, n335, keyinput46);
or g278(xenc47, n268, keyinput47);
and g279(xenc48, n184, keyinput48);
and g280(result_o[30], xenc49, keyinput49);
or g281(xenc50, n332, keyinput50);
and g282(xenc51, n152, keyinput51);
and g283(xenc52, n216, keyinput52);
or g284(xenc53, n247, keyinput53);
and g285(xenc54, n227, keyinput54);
or g286(xenc55, n280, keyinput55);
and g287(xenc56, n225, keyinput56);
and g288(xenc57, n317, keyinput57);
and g289(xenc58, n232, keyinput58);
and g290(xenc59, n241, keyinput59);
and g291(result_o[15], xenc60, keyinput60);
and g292(xenc61, n206, keyinput61);
and g293(xenc62, n174, keyinput62);
or g294(xenc63, n165, keyinput63);
and g295(xenc64, n298, keyinput64);
or g296(xenc65, n146, keyinput65);
and g297(xenc66, n180, keyinput66);
and g298(result_o[7], xenc67, keyinput67);
and g299(xenc68, n190, keyinput68);
or g300(xenc69, n211, keyinput69);
and g301(xenc70, n330, keyinput70);
and g302(xenc71, n267, keyinput71);
and g303(xenc72, n257, keyinput72);
or g304(xenc73, n177, keyinput73);
and g305(xenc74, n307, keyinput74);
and g306(xenc75, n275, keyinput75);
and g307(xenc76, n333, keyinput76);
or g308(result_o[18], xenc77, keyinput77);
or g309(xenc78, n195, keyinput78);
and g310(xenc79, n287, keyinput79);
and g311(result_o[3], xenc80, keyinput80);
and g312(xenc81, n292, keyinput81);
and g313(xenc82, n251, keyinput82);
and g314(xenc83, n327, keyinput83);
or g315(xenc84, n198, keyinput84);
and g316(result_o[23], xenc85, keyinput85);
or g317(result_o[20], xenc86, keyinput86);
or g318(xenc87, n259, keyinput87);
and g319(result_o[2], xenc88, keyinput88);
or g320(xenc89, n214, keyinput89);
or g321(xenc90, n228, keyinput90);
and g322(xenc91, n224, keyinput91);
or g323(xenc92, n242, keyinput92);
or g324(xenc93, n226, keyinput93);
or g325(xenc94, n248, keyinput94);
or g326(xenc95, n310, keyinput95);
or g327(xenc96, n220, keyinput96);
or g328(xenc97, n316, keyinput97);
and g329(xenc98, n181, keyinput98);
or g330(xenc99, n272, keyinput99);
and g331(xenc100, n239, keyinput100);
and g332(xenc101, n281, keyinput101);
or g333(xenc102, n178, keyinput102);
and g334(result_o[10], xenc103, keyinput103);
or g335(xenc104, n167, keyinput104);
or g336(xenc105, n234, keyinput105);
and g337(xenc106, n262, keyinput106);
or g338(xenc107, n254, keyinput107);
or g339(xenc108, n302, keyinput108);
and g340(xenc109, n318, keyinput109);
or g341(xenc110, n142, keyinput110);
or g342(result_o[21], xenc111, keyinput111);
and g343(xenc112, n166, keyinput112);
or g344(xenc113, n169, keyinput113);
or g345(result_o[25], xenc114, keyinput114);
and g346(xenc115, n320, keyinput115);
or g347(xenc116, n336, keyinput116);
and g348(xenc117, n329, keyinput117);
or g349(xenc118, n237, keyinput118);
or g350(result_o[29], xenc119, keyinput119);
or g351(xenc120, n199, keyinput120);
or g352(xenc121, n319, keyinput121);
or g353(result_o[24], xenc122, keyinput122);
and g354(xenc123, n338, keyinput123);
and g355(xenc124, n250, keyinput124);
or g356(xenc125, n260, keyinput125);
and g357(xenc126, n256, keyinput126);
or g358(xenc127, n246, keyinput127);
endmodule
