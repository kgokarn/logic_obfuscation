// Verilog File 
module broken_array_multiplier8_xor_enc64(op1_i,op2_i,keyinput,product_o);

input [7:0] op1_i,op2_i;
input [63:0] keyinput;

output [15:0] product_o;

wire n203, xenc15, xenc53, n205, n206, xenc12, n223, n238, n237, 
n230, n239, n229, n231, n236, n234, n258, n257, n256, n254, 
xenc45, n283, n281, n279, n269, n298, n275, xenc57, n326, n208, 
n327, n328, n325, n347, n348, n330, n349, xenc54, n355, n356, 
n319, n359, xenc35, n296, n301, n361, n307, xenc14, n310, n383, 
n384, n385, n386, xenc62, n391, n352, n392, n393, n390, n398, 
n399, n341, n402, n373, n372, n370, n441, n442, n443, n444, 
xenc19, n445, xenc31, n408, n461, xenc33, n429, n467, n468, n465, 
n417, n469, n409, n224, n225, n219, n221, n357, n358, n400, 
n401, n463, n464, n462, xenc52, n265, n276, n273, n297, xenc8, 
xenc48, n289, n293, n295, n333, xenc63, xenc60, n456, n436, n457, 
n458, n455, n250, n259, n248, n251, n290, n282, xenc2, n264, 
n334, n335, xenc20, n321, xenc30, n336, n291, xenc32, n294, n292, 
n260, n261, n263, n419, n420, n421, n284, xenc36, xenc26, n288, 
n286, n287, n285, n277, xenc42, n280, n278, n252, n253, n255, 
n374, n375, n313, n376, n449, n450, n430, n431, n451, n377, 
n378, n342, n343, n379, n246, n247, n249, n232, xenc40, n235, 
n233, n452, n453, n437, n438, n454, n422, n423, n424, n473, 
xenc25, n475, n474, n476, n477, xenc21, n478, n308, xenc22, xenc1, 
n309, n311, xenc37, n447, n446, n448, n302, n299, n267, n270, 
n415, xenc28, n244, n266, n242, n245, n351, n214, n353, n354, 
n329, xenc24, n212, n331, xenc51, n394, n395, n216, n396, n397, 
n435, xenc6, xenc41, n364, n366, n403, n318, n204, xenc13, n340, 
xenc11, n428, xenc5, n312, xenc23, n360, n315, n316, n317, n404, 
n405, xenc47, n407, n380, n381, xenc27, n382, xenc58, n338, n320, 
n337, n339, n368, xenc39, n306, n371, n369, n271, n272, xenc9, 
n274, xenc3, n388, n387, n389, n344, xenc49, xenc17, n345, n346, 
xenc61, n323, n209, xenc10, n322, xenc7, n324, n300, n432, xenc16, 
n434, n433, xenc43, n268, xenc46, n471, n470, n472, n314, n240, 
n241, n243, n226, n227, n228, n425, n426, n427, n362, xenc29, 
n365, n363, n413, xenc50, n412, xenc0, n414, n416, n303, xenc59, 
n305, n304, n207, xenc55, n222, n460, xenc38, n482, n481, n479, 
xenc18, n480, n220, n485, n486, n466, n459, n440, n483, n484, 
n439, n218, xenc56, n418, n410, n367, n202, n411, n350, n406, 
n210, n332, n262, n213, n211, xenc4, n215, xenc34, n487, xenc44;

xor g0(xenc53, n203, xenc15);
xor g1(n203, n205, n206);
xor g2(product_o[14], xenc12, n223);
xor g3(product_o[13], n238, n237);
xor g4(n237, n230, n239);
xor g5(n239, n229, n231);
xor g6(n238, n236, n234);
xor g7(product_o[12], n258, n257);
xor g8(n258, n256, n254);
xor g9(product_o[11], xenc45, n283);
xor g10(n283, n281, n279);
xor g11(n275, n269, n298);
xor g12(n208, xenc57, n326);
xor g13(n325, n327, n328);
xor g14(n330, n347, n348);
xor g15(n347, n349, xenc54);
xor g16(n319, n355, n356);
xor g17(n296, n359, xenc35);
xor g18(n307, n301, n361);
xor g19(n359, xenc14, n310);
xor g20(n348, n383, n384);
xor g21(n383, n385, n386);
xor g22(n352, xenc62, n391);
xor g23(n390, n392, n393);
xor g24(n341, n398, n399);
xor g25(n355, n402, n373);
xor g26(n402, n372, n370);
xor g27(n384, n441, n442);
xor g28(n442, n443, n444);
xor g29(n398, xenc19, n445);
xor g30(n445, xenc31, n408);
xor g31(n429, n461, xenc33);
xor g32(n465, n467, n468);
xor g33(n409, n417, n469);
nand g34(n219, n224, n225);
or g35(n221, n225, n224);
xnor g36(n356, n357, n358);
xnor g37(n399, n400, n401);
xnor g38(n462, n463, n464);
xnor g39(n265, xenc52, n275);
xnor g40(n297, n276, n273);
xnor g41(n289, xenc8, xenc48);
xnor g42(n333, n293, n295);
xnor g43(n441, n465, xenc63);
xnor g44(n436, xenc60, n456);
xnor g45(n455, n457, n458);
xnor g46(n257, n250, n259);
xnor g47(n259, n248, n251);
xnor g48(n282, n265, n290);
xnor g49(n290, xenc2, n264);
nand g50(n295, n334, n335);
or g51(n334, n319, xenc20);
nand g52(n335, n321, xenc30);
nand g53(n336, xenc20, n319);
nand g54(n264, n291, xenc32);
nand g55(n291, xenc8, n295);
nand g56(n292, n293, n294);
or g57(n294, n295, xenc8);
nand g58(n251, n260, n261);
nand g59(n260, n265, n264);
nand g60(n261, xenc2, n263);
or g61(n263, n264, n265);
nand g62(n372, n419, n420);
nand g63(n419, n398, n401);
nand g64(n420, n400, n421);
or g65(n421, n401, n398);
nand g66(n281, n284, xenc36);
nand g67(n284, xenc26, n288);
nand g68(n285, n286, n287);
or g69(n287, n288, xenc26);
nand g70(n256, n277, xenc42);
nand g71(n277, xenc45, n281);
nand g72(n278, n279, n280);
or g73(n280, n281, xenc45);
nand g74(n236, n252, n253);
nand g75(n252, n257, n256);
nand g76(n253, n254, n255);
or g77(n255, n256, n257);
nand g78(n313, n374, n375);
nand g79(n374, n355, n358);
nand g80(n375, n357, n376);
or g81(n376, n355, n358);
and g82(n444, n449, n450);
or g83(n449, n429, n430);
nand g84(n450, n431, n451);
nand g85(n451, n430, n429);
nand g86(n358, n377, n378);
or g87(n377, n341, n342);
nand g88(n378, n343, n379);
nand g89(n379, n342, n341);
and g90(n230, n246, n247);
nand g91(n246, n250, n251);
nand g92(n247, n248, n249);
or g93(n249, n250, n251);
nand g94(n225, n232, xenc40);
nand g95(n232, n237, n236);
nand g96(n233, n234, n235);
or g97(n235, n236, n237);
and g98(n430, n452, n453);
or g99(n452, n437, n438);
nand g100(n453, n436, n454);
nand g101(n454, n437, n438);
nand g102(n401, n422, n423);
nand g103(n422, n384, n385);
nand g104(n423, n386, n424);
or g105(n424, n385, n384);
nand g106(n468, n473, xenc25);
nand g107(n473, n461, n464);
nand g108(n474, n463, n475);
or g109(n475, n464, n461);
nand g110(n464, n476, n477);
nand g111(n476, n457, n456);
nand g112(n477, n458, xenc21);
or g113(n478, n456, n457);
and g114(n276, n308, xenc22);
nand g115(n308, xenc35, xenc14);
nand g116(n309, n310, xenc1);
or g117(n311, xenc35, xenc14);
and g118(n408, xenc37, n447);
or g119(n446, n441, n444);
nand g120(n447, n443, n448);
nand g121(n448, n444, n441);
xnor g122(n361, n302, n299);
xnor g123(n298, n267, n270);
xnor g124(n469, n415, xenc28);
xnor g125(n250, n244, n266);
xnor g126(n266, n242, n245);
xnor g127(n214, n351, n352);
xnor g128(n351, n353, n354);
xnor g129(n212, n329, xenc24);
xnor g130(n329, n331, xenc51);
xnor g131(n216, n394, n395);
xnor g132(n394, n396, n397);
xnor g133(n395, n435, n436);
xnor g134(n435, n437, n438);
xnor g135(n373, xenc6, xenc41);
xnor g136(n403, n364, n366);
xnor g137(n204, n318, n319);
xnor g138(n318, xenc20, n321);
xnor g139(n326, xenc13, n341);
xnor g140(n340, n342, n343);
xnor g141(n391, xenc11, n429);
xnor g142(n428, n430, n431);
xnor g143(n312, xenc5, n307);
xnor g144(n360, xenc23, n267);
nand g145(n288, n315, n316);
nand g146(n315, n206, n205);
nand g147(n316, xenc15, n317);
or g148(n317, n205, n206);
nand g149(n366, n404, n405);
or g150(n404, xenc19, n408);
nand g151(n405, xenc31, xenc47);
nand g152(n407, n408, xenc19);
and g153(n342, n380, n381);
nand g154(n380, xenc54, n349);
nand g155(n381, n348, xenc27);
or g156(n382, n349, xenc54);
and g157(n320, xenc58, n338);
nand g158(n337, n328, n327);
nand g159(n338, n326, n339);
or g160(n339, n327, n328);
and g161(n306, n368, xenc39);
nand g162(n368, n373, n372);
nand g163(n369, n370, n371);
or g164(n371, n372, n373);
and g165(n244, n271, n272);
or g166(n271, n275, n276);
nand g167(n272, n273, xenc9);
nand g168(n274, n275, n276);
nand g169(n349, xenc3, n388);
or g170(n387, n353, n354);
nand g171(n388, n352, n389);
nand g172(n389, n353, n354);
nand g173(n327, n344, xenc49);
nand g174(n344, n331, xenc51);
nand g175(n345, xenc24, xenc17);
or g176(n346, n331, xenc51);
nand g177(n205, xenc61, n323);
or g178(n322, n209, xenc10);
nand g179(n323, xenc7, n324);
nand g180(n324, n209, xenc10);
nand g181(n270, n299, n300);
nand g182(n300, n301, n302);
nand g183(n392, n432, xenc16);
or g184(n432, n396, n397);
nand g185(n433, n395, n434);
nand g186(n434, n396, n397);
and g187(n242, n267, xenc43);
nand g188(n268, n269, n270);
and g189(n417, xenc46, n471);
nand g190(n470, xenc63, n468);
nand g191(n471, n467, n472);
or g192(n472, n468, xenc63);
xnor g193(product_o[10], xenc26, n314);
xnor g194(n314, n286, n288);
nand g195(n229, n240, n241);
or g196(n240, n245, n244);
nand g197(n241, n242, n243);
nand g198(n243, n244, n245);
nand g199(n224, n226, n227);
or g200(n226, n231, n230);
nand g201(n227, n228, n229);
nand g202(n228, n230, n231);
nand g203(n385, n425, n426);
nand g204(n425, n393, n392);
nand g205(n426, n391, n427);
or g206(n427, n392, n393);
and g207(n301, n362, xenc29);
nand g208(n362, xenc6, n366);
nand g209(n363, n364, n365);
or g210(n365, n366, xenc6);
nand g211(n412, n413, xenc50);
or g212(n413, xenc28, n417);
nand g213(n414, n415, xenc0);
nand g214(n416, n417, xenc28);
and g215(n269, n303, xenc59);
or g216(n303, n307, xenc23);
nand g217(n304, n267, n305);
nand g218(n305, xenc23, n307);
xnor g219(product_o[8], n207, xenc7);
xnor g220(n207, n209, xenc10);
nand g221(n223, op2_i[7], op1_i[7]);
nand g222(n222, xenc55, n219);
and g223(n457, op2_i[2], n460, op1_i[2]);
xnor g224(n460, xenc38, n482);
nand g225(n481, op1_i[3], op2_i[1]);
and g226(n482, op1_i[4], op2_i[0]);
xnor g227(n456, n479, xenc18);
nand g228(n479, op1_i[4], op2_i[1]);
and g229(n480, op1_i[5], op2_i[0]);
nand g230(product_o[15], n219, n220);
nand g231(n220, op1_i[7], xenc55, op2_i[7]);
xnor g232(n466, n485, n486);
nand g233(n485, op1_i[6], op2_i[1]);
and g234(n486, op1_i[7], op2_i[0]);
xnor g235(n440, n459, n460);
nand g236(n459, op1_i[2], op2_i[2]);
xnor g237(n461, n483, n484);
nand g238(n483, op1_i[5], op2_i[1]);
and g239(n484, op1_i[6], op2_i[0]);
xnor g240(n218, n439, n440);
nand g241(n439, op1_i[1], op2_i[3]);
nand g242(n209, op1_i[0], xenc56, op2_i[7]);
nand g243(n353, op1_i[0], n216, op2_i[5]);
nand g244(n437, op2_i[3], n440, op1_i[1]);
nand g245(n396, op2_i[4], n218, op1_i[0]);
nand g246(n418, op2_i[2], op1_i[6]);
nand g247(n438, op2_i[3], op1_i[2]);
nand g248(n397, op2_i[4], op1_i[1]);
nand g249(n354, op2_i[5], op1_i[1]);
nand g250(n302, op1_i[7], n412);
and g251(n367, n302, n410);
nand g252(n410, n202, n411);
nand g253(n411, op2_i[2], op1_i[7]);
not g254(n202, n412);
and g255(n458, op1_i[3], op2_i[2]);
and g256(n431, op2_i[3], op1_i[3]);
and g257(n393, op2_i[4], op1_i[2]);
and g258(n350, op2_i[5], op1_i[2]);
and g259(n463, op1_i[4], op2_i[2]);
and g260(n415, op2_i[1], op1_i[7]);
and g261(n400, op2_i[4], op1_i[4]);
and g262(n364, op2_i[3], op1_i[6]);
and g263(n331, op2_i[6], op1_i[0], n214);
and g264(n386, op2_i[4], op1_i[3]);
and g265(n467, op1_i[5], op2_i[2]);
and g266(n443, op2_i[3], op1_i[4]);
and g267(n406, op2_i[3], op1_i[5]);
and g268(n267, op2_i[4], op1_i[6]);
nand g269(n245, op2_i[5], op1_i[7]);
nand g270(n210, op2_i[7], op1_i[1]);
and g271(n332, op2_i[6], op1_i[1]);
and g272(n343, op2_i[5], op1_i[3]);
and g273(n299, op2_i[3], op1_i[7]);
and g274(n321, op2_i[6], op1_i[3]);
and g275(n273, op2_i[5], op1_i[6]);
and g276(n328, op2_i[6], op1_i[2]);
and g277(n206, op2_i[7], op1_i[2]);
and g278(n357, op2_i[5], op1_i[4]);
and g279(n293, op2_i[6], op1_i[4]);
and g280(n286, op2_i[7], op1_i[3]);
and g281(n262, op2_i[6], op1_i[5]);
and g282(n248, op2_i[6], op1_i[6]);
xnor g283(product_o[6], n213, n214);
nand g284(n213, op2_i[6], op1_i[0]);
xnor g285(xenc4, n211, xenc56);
nand g286(n211, op2_i[7], op1_i[0]);
and g287(n370, op2_i[4], op1_i[5]);
and g288(n310, op2_i[5], op1_i[5]);
xnor g289(xenc34, n215, n216);
nand g290(n215, op2_i[5], op1_i[0]);
nand g291(n231, op2_i[6], op1_i[7]);
xnor g292(product_o[4], n487, n218);
nand g293(n487, op2_i[4], op1_i[0]);
and g294(n279, op2_i[7], op1_i[4]);
and g295(n254, op2_i[7], op1_i[5]);
and g296(n234, op2_i[7], op1_i[6]);
and g297(product_o[0], op2_i[0], op1_i[0]);
and g298(product_o[1], op2_i[1], op1_i[0]);
and g299(product_o[2], op2_i[2], op1_i[0]);
and g300(xenc44, op2_i[3], op1_i[0]);
xnor g301(xenc0, n416, keyinput[0]);
xnor g302(xenc1, n311, keyinput[1]);
xnor g303(xenc2, n262, keyinput[2]);
xor g304(xenc3, n387, keyinput[3]);
xor g305(product_o[7], xenc4, keyinput[4]);
xnor g306(xenc5, n360, keyinput[5]);
xor g307(xenc6, n367, keyinput[6]);
xor g308(xenc7, n208, keyinput[7]);
xnor g309(xenc8, n296, keyinput[8]);
xnor g310(xenc9, n274, keyinput[9]);
xor g311(xenc10, n210, keyinput[10]);
xor g312(xenc11, n428, keyinput[11]);
xnor g313(xenc12, n222, keyinput[12]);
xnor g314(xenc13, n340, keyinput[13]);
xor g315(xenc14, n313, keyinput[14]);
xnor g316(xenc15, n204, keyinput[15]);
xor g317(xenc16, n433, keyinput[16]);
xor g318(xenc17, n346, keyinput[17]);
xor g319(xenc18, n480, keyinput[18]);
xnor g320(xenc19, n409, keyinput[19]);
xor g321(xenc20, n320, keyinput[20]);
xor g322(xenc21, n478, keyinput[21]);
xnor g323(xenc22, n309, keyinput[22]);
xor g324(xenc23, n306, keyinput[23]);
xnor g325(xenc24, n330, keyinput[24]);
xnor g326(xenc25, n474, keyinput[25]);
xnor g327(xenc26, n289, keyinput[26]);
xnor g328(xenc27, n382, keyinput[27]);
xor g329(xenc28, n418, keyinput[28]);
xnor g330(xenc29, n363, keyinput[29]);
xor g331(xenc30, n336, keyinput[30]);
xor g332(xenc31, n406, keyinput[31]);
xnor g333(xenc32, n292, keyinput[32]);
xor g334(xenc33, n462, keyinput[33]);
xnor g335(product_o[5], xenc34, keyinput[34]);
xor g336(xenc35, n312, keyinput[35]);
xor g337(xenc36, n285, keyinput[36]);
xnor g338(xenc37, n446, keyinput[37]);
xor g339(xenc38, n481, keyinput[38]);
xor g340(xenc39, n369, keyinput[39]);
xnor g341(xenc40, n233, keyinput[40]);
xnor g342(xenc41, n403, keyinput[41]);
xnor g343(xenc42, n278, keyinput[42]);
xor g344(xenc43, n268, keyinput[43]);
xnor g345(product_o[3], xenc44, keyinput[44]);
xnor g346(xenc45, n282, keyinput[45]);
xor g347(xenc46, n470, keyinput[46]);
xor g348(xenc47, n407, keyinput[47]);
xor g349(xenc48, n333, keyinput[48]);
xor g350(xenc49, n345, keyinput[49]);
xnor g351(xenc50, n414, keyinput[50]);
xor g352(xenc51, n332, keyinput[51]);
xnor g353(xenc52, n297, keyinput[52]);
xnor g354(product_o[9], xenc53, keyinput[53]);
xnor g355(xenc54, n350, keyinput[54]);
xor g356(xenc55, n221, keyinput[55]);
xor g357(xenc56, n212, keyinput[56]);
xnor g358(xenc57, n325, keyinput[57]);
xor g359(xenc58, n337, keyinput[58]);
xnor g360(xenc59, n304, keyinput[59]);
xnor g361(xenc60, n455, keyinput[60]);
xnor g362(xenc61, n322, keyinput[61]);
xor g363(xenc62, n390, keyinput[62]);
xor g364(xenc63, n466, keyinput[63]);
endmodule
