// Verilog File 
module ripple_carry_adder32_xor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n886, xenc96, n812, xenc30, xenc25, xenc117, xenc120, xenc47, xenc119, 
n820, xenc70, xenc104, xenc64, xenc93, xenc41, xenc35, n857, n859, n863, 
n864, xenc81, xenc126, xenc94, n871, xenc123, n875, xenc105, xenc10, xenc71, 
n887, xenc127, n894, n895, xenc6, n907, xenc68, xenc121, xenc62, n913, 
n921, xenc33, n927, xenc42, xenc45, xenc114, n837, xenc28, xenc108, n841, 
xenc54, n915, xenc72, n911, xenc74, n998, n995, n931, n977, n965, 
n959, xenc80, n957, n996, n800, n900, n901, n893, xenc84, n974, 
xenc21, n966, n946, xenc85, n948, n985, xenc52, n1000, n865, n967, 
xenc12, n969, n976, xenc77, n830, n827, n937, n943, n938, n922, 
xenc43, n855, xenc87, n981, xenc59, n840, n983, n968, n818, xenc24, 
n904, n903, xenc36, n799, n896, xenc46, n880, n823, xenc22, n849, 
xenc91, n848, n1003, xenc97, n970, n897, xenc4, n910, n971, xenc29, 
xenc40, n972, xenc50, n973, xenc89, n925, xenc57, xenc39, n975, xenc125, 
n942, n815, n816, n892, xenc15, n890, xenc118, n978, n979, n990, 
n980, n991, n982, n836, xenc26, n984, xenc99, n987, n986, n988, 
xenc116, n989, xenc109, n797, xenc19, n916, n845, xenc58, n992, n993, 
n933, n801, n934, n994, n831, n997, n999, xenc7, n862, xenc65, 
n1001, n1002, xenc37, n1005, n1004, n930, xenc110, xenc83, n1006, n1007, 
xenc8, n884, n824, n1012, n1011, xenc103, n834, n835, n833, xenc17, 
n850, n852, xenc9, n853, n851, xenc86, xenc60, xenc5, n1008, xenc106, 
n832, n1009, n802, xenc23, n939, n944, n940, xenc82, n945, n803, 
n898, n917, xenc49, xenc75, n798, n1010, xenc18, n814, n808, xenc53, 
xenc56, xenc95, n889, n885, xenc124, xenc31, n867, xenc107, xenc11, n902, 
n879, xenc44, xenc32, n924, xenc100, xenc3, xenc79, n861, n947, xenc78, 
xenc66, xenc101, n956, xenc48, n914, n846, xenc34, n826, n817, n958, 
n955, n954, n952, n847, n873, n919, xenc27, n912, n962, xenc73, 
n960, n963, n877, xenc51, n876, xenc13, n821, xenc102, n928, n810, 
xenc0, xenc63, xenc1, xenc88, xenc55, n868, n869, xenc98, n905, n953, 
xenc115, n951, n819, xenc112, n828, n839, xenc69, n888, n891, n920, 
n918, n935, n811, xenc67, n858, n856, n854, n874, n872, n878, 
xenc14, n926, n809, xenc113, xenc122, xenc20, n860, xenc76, xenc61, n881, 
n883, xenc111, n906, n923, xenc2, n932, n936, n961, n822, xenc92, 
n825, n796, n866, n870, n882, n909, n929, xenc38, xenc90, xenc16, 
n941;

or g0(n886, add2_i[0], add1_i[0]);
xor g1(xenc30, xenc96, n812);
xor g2(xenc117, add2_i[6], xenc25);
xor g3(xenc47, add2_i[5], xenc120);
xor g4(result_o[3], xenc119, n820);
xor g5(n820, add2_i[3], add1_i[3]);
xor g6(xenc104, xenc70, add2_i[2]);
xor g7(xenc93, add2_i[28], xenc64);
xor g8(result_o[27], add2_i[27], xenc41);
xor g9(result_o[26], xenc35, n857);
xor g10(result_o[25], n859, add2_i[25]);
xor g11(xenc81, n863, n864);
xor g12(n864, add2_i[24], add1_i[24]);
xor g13(xenc94, add2_i[23], xenc126);
xor g14(xenc123, add2_i[22], n871);
xor g15(xenc105, add2_i[21], n875);
xor g16(result_o[1], xenc10, xenc71);
xor g17(n887, add2_i[1], add1_i[1]);
xor g18(result_o[19], xenc127, add2_i[19]);
xor g19(xenc6, n894, n895);
xor g20(result_o[15], add2_i[15], n907);
xor g21(xenc62, xenc68, xenc121);
xor g22(n913, add2_i[14], add1_i[14]);
xor g23(result_o[12], n921, add2_i[12]);
xor g24(xenc42, xenc33, n927);
xor g25(n927, add2_i[11], add1_i[11]);
xor g26(result_o[10], xenc45, add2_i[10]);
xor g27(n837, xenc114, add1_i[2]);
nand g28(n841, xenc28, xenc108);
nand g29(n911, xenc54, n915, xenc72);
nand g30(n995, xenc74, add2_i[28], add1_i[29], n998);
xor g31(n977, n931, add1_i[10]);
nand g32(n957, n965, n959, xenc80);
not g33(n965, add1_i[3]);
nand g34(n996, n841, add1_i[28], add1_i[29]);
nand g35(n893, n800, n900, n901);
nor g36(n974, xenc84, add1_i[11]);
not g37(n966, xenc21);
and g38(n985, n946, xenc85, n948);
nor g39(n1000, xenc52, add1_i[24]);
not g40(n967, n865);
nand g41(n969, xenc12, add2_i[16], add1_i[17]);
nand g42(n827, n976, xenc77, n996, n830);
nand g43(n938, n937, n943, add2_i[6]);
xor g44(n921, n922, add1_i[12]);
xor g45(n871, xenc43, add1_i[22]);
xor g46(n859, n855, add1_i[25]);
nor g47(n840, xenc87, n981, xenc59);
not g48(n968, n983);
xnor g49(result_o[0], add2_i[0], add1_i[0]);
xor g50(xenc24, add2_i[4], n818);
xnor g51(n903, n904, add1_i[16]);
and g52(n896, add2_i[17], xenc36, n799);
xnor g53(n880, xenc46, add1_i[20]);
xor g54(xenc22, n823, add2_i[31]);
and g55(n848, n849, xenc91);
not g56(n1003, add1_i[4]);
nand g57(n897, xenc97, n970);
or g58(n970, n800, n901);
nand g59(n971, xenc4, n910);
nand g60(n972, xenc29, xenc40);
nand g61(n973, xenc50, add2_i[10]);
nand g62(n925, n973, xenc89);
nand g63(n975, xenc57, xenc39);
not g64(n976, add1_i[30]);
and g65(n815, xenc125, n942);
and g66(n816, n943, n937);
nand g67(n890, n892, xenc15);
nor g68(n978, xenc118, add1_i[18]);
and g69(n979, xenc120, xenc85);
nor g70(n998, xenc59, n981);
and g71(n980, add1_i[28], n990);
and g72(n981, n991, add1_i[28]);
or g73(n982, n991, add1_i[28], n990);
or g74(n983, n991, add1_i[28], n990);
or g75(n836, n991, add1_i[28], n990);
nor g76(n984, n979, xenc26);
nor g77(n937, xenc99, xenc26);
nor g78(n986, n987, n946);
not g79(n987, add1_i[6]);
and g80(n988, add2_i[5], add1_i[6]);
or g81(n989, xenc116, add1_i[13]);
nor g82(n990, xenc108, xenc109);
nor g83(n991, n797, xenc19);
or g84(n916, xenc116, add1_i[13]);
nor g85(n845, n797, xenc19);
nand g86(n992, add2_i[27], xenc58);
nand g87(n993, xenc4, n910);
nand g88(n994, n933, n801, n934);
and g89(n831, xenc77, n996);
not g90(n997, add1_i[29]);
nand g91(n999, xenc126, add2_i[23]);
nand g92(n862, n999, xenc7);
nand g93(n1001, xenc65, add2_i[13]);
not g94(n1002, add1_i[14]);
xnor g95(n818, xenc37, n1003);
not g96(n1005, add1_i[21]);
not g97(n1004, add1_i[10]);
xnor g98(n930, n931, n1004);
xnor g99(n875, xenc110, xenc83);
not g100(n1006, add1_i[19]);
not g101(n1007, add1_i[31]);
xnor g102(n884, xenc8, n1006);
xnor g103(n823, n824, n1007);
not g104(n1012, add1_i[15]);
not g105(n1011, add1_i[23]);
nand g106(n830, xenc103, add2_i[29]);
nand g107(n833, n834, n997, n835);
nand g108(n850, add2_i[26], xenc17);
nand g109(n851, n852, xenc9, n853);
not g110(n801, add1_i[9]);
xnor g111(n857, add2_i[26], xenc9);
or g112(n948, xenc86, add1_i[5]);
xor g113(result_o[30], xenc60, xenc5);
xor g114(n1008, add1_i[30], add2_i[30]);
xor g115(result_o[29], xenc106, n832);
xor g116(n1009, add1_i[29], add2_i[29]);
nand g117(n834, add1_i[28], n841);
not g118(n802, add1_i[8]);
xnor g119(result_o[20], add2_i[20], xenc23);
nand g120(n933, add2_i[8], n939);
nand g121(n940, add2_i[7], n944);
nand g122(n852, add2_i[25], xenc82);
nand g123(n945, add2_i[6], n943);
not g124(n803, add1_i[7]);
xnor g125(n894, add1_i[18], add2_i[18]);
xnor g126(result_o[17], add2_i[17], n898);
xnor g127(xenc49, add2_i[13], n917);
xnor g128(result_o[16], add2_i[16], n903);
not g129(n800, add1_i[17]);
xnor g130(n812, add2_i[8], xenc75);
not g131(n798, add1_i[26]);
xnor g132(xenc18, add2_i[7], n1010);
nand g133(n1010, n814, xenc29);
xnor g134(xenc53, add2_i[9], n808);
not g135(n797, add1_i[27]);
nand g136(n943, n946, n987, xenc56);
nand g137(n885, xenc95, n889);
xnor g138(n867, xenc124, xenc31);
xnor g139(n907, xenc107, xenc11);
or g140(n902, n904, add1_i[16]);
or g141(n879, xenc46, add1_i[20]);
nand g142(n917, n915, xenc65);
nand g143(n910, xenc44, add2_i[14]);
nand g144(n924, xenc32, add2_i[11]);
nand g145(n922, xenc100, xenc3);
nand g146(n855, xenc57, xenc39);
nand g147(n861, add2_i[24], xenc79);
nand g148(n947, n948, add2_i[5]);
nand g149(n824, xenc78, xenc66);
nand g150(n956, xenc101, add2_i[3]);
nand g151(n914, xenc48, add2_i[13]);
and g152(n846, xenc28, xenc58);
nand g153(n826, xenc34, add2_i[30]);
and g154(n817, n946, n948);
nand g155(n958, add1_i[2], xenc114);
nand g156(n954, n956, n955);
nand g157(n952, add1_i[4], xenc37);
nand g158(n847, xenc19, n797);
nand g159(n873, add1_i[21], xenc110);
nand g160(n889, n890, add2_i[18]);
nand g161(n919, add1_i[12], n922);
nand g162(n912, xenc27, n915);
nand g163(n900, xenc12, add2_i[16]);
nand g164(n960, n962, xenc73);
nand g165(n962, n963, add2_i[1]);
nand g166(n876, n877, xenc51);
nand g167(n877, xenc13, add2_i[20]);
nand g168(n821, add1_i[31], n824);
nand g169(n863, n865, xenc102);
nand g170(n865, xenc124, add1_i[23]);
nand g171(n928, n931, add1_i[10]);
nand g172(n931, n810, xenc0);
nand g173(n939, xenc63, xenc75, xenc29);
nand g174(n946, add1_i[5], xenc86);
nand g175(n832, n834, xenc1);
nand g176(n868, xenc88, xenc55);
nand g177(n869, xenc43, add1_i[22]);
nand g178(n905, xenc98, add1_i[15]);
nand g179(n915, add1_i[13], xenc116);
nand g180(n951, n953, xenc115);
nand g181(n819, n959, xenc80);
nand g182(n828, xenc112, n830);
nand g183(n839, add2_i[28], xenc64);
nand g184(n849, add1_i[26], xenc35);
nand g185(n888, add1_i[18], xenc69);
nand g186(n891, n892, n799);
nand g187(n918, n919, n920);
nand g188(n810, n935, add1_i[9]);
nand g189(n934, add1_i[8], n811);
nand g190(n898, xenc36, n799);
nand g191(n835, add2_i[28], xenc67);
nand g192(n856, n853, n858);
nand g193(n853, add1_i[25], n975);
or g194(n854, n975, add1_i[25]);
nand g195(n872, n874, n873);
nand g196(n878, add1_i[20], xenc46);
nand g197(n892, add2_i[17], xenc36);
nand g198(n926, xenc21, xenc14);
nand g199(n935, n933, n934);
nand g200(n809, n933, n801, n934);
nand g201(n811, xenc29, xenc40);
nand g202(result_o[32], xenc113, xenc122);
nand g203(n808, xenc20, n810);
nand g204(n860, add1_i[24], n863);
nand g205(n881, xenc76, xenc61);
nand g206(n883, add2_i[19], xenc127);
nand g207(n901, add1_i[16], n904);
nand g208(n904, xenc111, n906);
nand g209(n923, add1_i[11], xenc33);
nand g210(n932, add2_i[9], xenc2);
nand g211(n936, add2_i[7], n814);
nand g212(n955, add1_i[3], xenc119);
nand g213(n961, add1_i[1], xenc10);
or g214(n963, xenc10, add1_i[1]);
nand g215(n822, add2_i[31], n823);
nor g216(n895, xenc92, xenc118);
nand g217(n825, add1_i[30], xenc5);
not g218(n796, n991);
nand g219(n858, n859, add2_i[25]);
nand g220(n866, add2_i[23], xenc126);
nand g221(n870, add2_i[22], n871);
nand g222(n874, add2_i[21], n875);
nand g223(n882, xenc8, add1_i[19]);
not g224(n799, xenc118);
nand g225(n906, add2_i[15], n907);
nand g226(n909, add1_i[14], xenc68);
nand g227(n920, add2_i[12], n921);
nand g228(n929, add2_i[10], xenc45);
nand g229(n944, xenc38, n803, xenc90);
nand g230(n814, xenc38, n803, xenc16);
nand g231(n942, add1_i[7], xenc25, add2_i[6]);
or g232(n941, xenc38, n803);
nand g233(n953, n818, add2_i[4]);
nand g234(n959, add2_i[2], xenc70);
xnor g235(xenc0, n932, keyinput0);
xor g236(xenc1, n839, keyinput1);
xnor g237(xenc2, n809, keyinput2);
xnor g238(xenc3, n923, keyinput3);
xnor g239(xenc4, n909, keyinput4);
xor g240(xenc5, n828, keyinput5);
xnor g241(result_o[18], xenc6, keyinput6);
xnor g242(xenc7, n1000, keyinput7);
xnor g243(xenc8, n885, keyinput8);
xnor g244(xenc9, n798, keyinput9);
xor g245(xenc10, n886, keyinput10);
xnor g246(xenc11, n1012, keyinput11);
xor g247(xenc12, n902, keyinput12);
xor g248(xenc13, n879, keyinput13);
xor g249(xenc14, n929, keyinput14);
xnor g250(xenc15, n978, keyinput15);
xor g251(xenc16, n938, keyinput16);
xnor g252(xenc17, n851, keyinput17);
xnor g253(result_o[7], xenc18, keyinput18);
xor g254(xenc19, n848, keyinput19);
xor g255(xenc20, n994, keyinput20);
xnor g256(xenc21, n928, keyinput21);
xnor g257(result_o[31], xenc22, keyinput22);
xor g258(xenc23, n880, keyinput23);
xnor g259(result_o[4], xenc24, keyinput24);
xor g260(xenc25, n816, keyinput25);
xnor g261(xenc26, n986, keyinput26);
xnor g262(xenc27, n914, keyinput27);
xor g263(xenc28, n796, keyinput28);
xnor g264(xenc29, n815, keyinput29);
xnor g265(result_o[8], xenc30, keyinput30);
xor g266(xenc31, n1011, keyinput31);
xnor g267(xenc32, n925, keyinput32);
xor g268(xenc33, n926, keyinput33);
xor g269(xenc34, n827, keyinput34);
xnor g270(xenc35, n856, keyinput35);
xnor g271(xenc36, n893, keyinput36);
xor g272(xenc37, n954, keyinput37);
xnor g273(xenc38, n984, keyinput38);
xor g274(xenc39, n860, keyinput39);
xor g275(xenc40, n936, keyinput40);
xor g276(xenc41, n846, keyinput41);
xor g277(result_o[11], xenc42, keyinput42);
xor g278(xenc43, n872, keyinput43);
xor g279(xenc44, n911, keyinput44);
xnor g280(xenc45, n930, keyinput45);
xor g281(xenc46, n881, keyinput46);
xnor g282(result_o[5], xenc47, keyinput47);
xnor g283(xenc48, n916, keyinput48);
xor g284(result_o[13], xenc49, keyinput49);
xnor g285(xenc50, n977, keyinput50);
xor g286(xenc51, n878, keyinput51);
xnor g287(xenc52, n967, keyinput52);
xnor g288(result_o[9], xenc53, keyinput53);
xnor g289(xenc54, n1002, keyinput54);
xnor g290(xenc55, n869, keyinput55);
xnor g291(xenc56, n947, keyinput56);
xnor g292(xenc57, n861, keyinput57);
xnor g293(xenc58, n847, keyinput58);
xor g294(xenc59, n980, keyinput59);
xor g295(xenc60, n1008, keyinput60);
xor g296(xenc61, n882, keyinput61);
xnor g297(result_o[14], xenc62, keyinput62);
xor g298(xenc63, n940, keyinput63);
xnor g299(xenc64, n840, keyinput64);
xnor g300(xenc65, n989, keyinput65);
xor g301(xenc66, n826, keyinput66);
xnor g302(xenc67, n982, keyinput67);
xor g303(xenc68, n912, keyinput68);
xor g304(xenc69, n891, keyinput69);
xor g305(xenc70, n837, keyinput70);
xor g306(xenc71, n887, keyinput71);
xnor g307(xenc72, n1001, keyinput72);
xor g308(xenc73, n961, keyinput73);
xnor g309(xenc74, n836, keyinput74);
xor g310(xenc75, n802, keyinput75);
xor g311(xenc76, n883, keyinput76);
xor g312(xenc77, n995, keyinput77);
xnor g313(xenc78, n825, keyinput78);
xnor g314(xenc79, n862, keyinput79);
xnor g315(xenc80, n958, keyinput80);
xnor g316(result_o[24], xenc81, keyinput81);
xor g317(xenc82, n854, keyinput82);
xnor g318(xenc83, n1005, keyinput83);
xnor g319(xenc84, n966, keyinput84);
xnor g320(xenc85, n988, keyinput85);
xnor g321(xenc86, n951, keyinput86);
xnor g322(xenc87, n968, keyinput87);
xnor g323(xenc88, n870, keyinput88);
xor g324(xenc89, n974, keyinput89);
xor g325(xenc90, n945, keyinput90);
xor g326(xenc91, n850, keyinput91);
xnor g327(xenc92, n896, keyinput92);
xnor g328(result_o[28], xenc93, keyinput93);
xnor g329(result_o[23], xenc94, keyinput94);
xnor g330(xenc95, n888, keyinput95);
xnor g331(xenc96, n972, keyinput96);
xor g332(xenc97, n969, keyinput97);
xnor g333(xenc98, n971, keyinput98);
xor g334(xenc99, n985, keyinput99);
xnor g335(xenc100, n924, keyinput100);
xnor g336(xenc101, n957, keyinput101);
xnor g337(xenc102, n866, keyinput102);
xor g338(xenc103, n833, keyinput103);
xor g339(result_o[2], xenc104, keyinput104);
xnor g340(result_o[21], xenc105, keyinput105);
xnor g341(xenc106, n1009, keyinput106);
xnor g342(xenc107, n993, keyinput107);
xor g343(xenc108, n992, keyinput108);
xnor g344(xenc109, n845, keyinput109);
xnor g345(xenc110, n876, keyinput110);
xnor g346(xenc111, n905, keyinput111);
xnor g347(xenc112, n831, keyinput112);
xnor g348(xenc113, n821, keyinput113);
xnor g349(xenc114, n960, keyinput114);
xor g350(xenc115, n952, keyinput115);
xnor g351(xenc116, n918, keyinput116);
xor g352(result_o[6], xenc117, keyinput117);
xor g353(xenc118, n897, keyinput118);
xnor g354(xenc119, n819, keyinput119);
xnor g355(xenc120, n817, keyinput120);
xor g356(xenc121, n913, keyinput121);
xnor g357(xenc122, n822, keyinput122);
xnor g358(result_o[22], xenc123, keyinput123);
xor g359(xenc124, n868, keyinput124);
xnor g360(xenc125, n941, keyinput125);
xnor g361(xenc126, n867, keyinput126);
xor g362(xenc127, n884, keyinput127);
endmodule
