module lower_part_or_carry_lookahead_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147;

  xor U119 ( result_o[9], n28, n29);
  xor U120 ( n29, add2_i[9], add1_i[9]);
  xor U121 ( result_o[8], n30, n31);
  xor U122 ( n31, add2_i[8], add1_i[8]);
  xor U123 ( result_o[31], n35, n36);
  xor U124 ( n36, add2_i[31], add1_i[31]);
  xor U125 ( result_o[30], n40, n41);
  xor U126 ( n41, add2_i[30], add1_i[30]);
  xor U127 ( result_o[29], n45, n46);
  xor U128 ( n46, add2_i[29], add1_i[29]);
  xor U129 ( result_o[28], n50, n51);
  xor U130 ( n51, add2_i[28], add1_i[28]);
  xor U131 ( result_o[27], n55, n56);
  xor U132 ( n56, add2_i[27], add1_i[27]);
  xor U133 ( result_o[26], n60, n61);
  xor U134 ( n61, add2_i[26], add1_i[26]);
  xor U135 ( result_o[25], n65, n66);
  xor U136 ( n66, add2_i[25], add1_i[25]);
  xor U137 ( result_o[24], n70, n71);
  xor U138 ( n71, add2_i[24], add1_i[24]);
  xor U139 ( result_o[23], n75, n76);
  xor U140 ( n76, add2_i[23], add1_i[23]);
  xor U141 ( result_o[22], n80, n81);
  xor U142 ( n81, add2_i[22], add1_i[22]);
  xor U143 ( result_o[21], n85, n86);
  xor U144 ( n86, add2_i[21], add1_i[21]);
  xor U145 ( result_o[20], n90, n91);
  xor U146 ( n91, add2_i[20], add1_i[20]);
  xor U147 ( result_o[19], n95, n96);
  xor U148 ( n96, add2_i[19], add1_i[19]);
  xor U149 ( result_o[18], n100, n101);
  xor U150 ( n101, add2_i[18], add1_i[18]);
  xor U151 ( result_o[17], n105, n106);
  xor U152 ( n106, add2_i[17], add1_i[17]);
  xor U153 ( result_o[16], n110, n111);
  xor U154 ( n111, add2_i[16], add1_i[16]);
  xor U155 ( result_o[15], n115, n116);
  xor U156 ( n116, add2_i[15], add1_i[15]);
  xor U157 ( result_o[14], n120, n121);
  xor U158 ( n121, add2_i[14], add1_i[14]);
  xor U159 ( result_o[13], n125, n126);
  xor U160 ( n126, add2_i[13], add1_i[13]);
  xor U161 ( result_o[12], n130, n131);
  xor U162 ( n131, add2_i[12], add1_i[12]);
  xor U163 ( result_o[11], n135, n136);
  xor U164 ( n136, add2_i[11], add1_i[11]);
  xor U165 ( result_o[10], n140, n141);
  xor U166 ( n141, add2_i[10], add1_i[10]);
  nand U167 ( result_o[7], n27, n26);
  nand U168 ( n28, n145, n146);
  nand U169 ( n145, add2_i[8], add1_i[8]);
  nand U170 ( n146, add1_i[7], n147, add2_i[7]);
  or U171 ( n147, add2_i[8], add1_i[8]);
  nand U172 ( n140, n142, n143);
  nand U173 ( n142, add1_i[9], n28);
  nand U174 ( n143, add2_i[9], n144);
  or U175 ( n144, n28, add1_i[9]);
  nand U176 ( n135, n137, n138);
  nand U177 ( n137, add1_i[10], n140);
  nand U178 ( n138, add2_i[10], n139);
  or U179 ( n139, n140, add1_i[10]);
  nand U180 ( n130, n132, n133);
  nand U181 ( n132, add1_i[11], n135);
  nand U182 ( n133, add2_i[11], n134);
  or U183 ( n134, n135, add1_i[11]);
  nand U184 ( n125, n127, n128);
  nand U185 ( n127, add1_i[12], n130);
  nand U186 ( n128, add2_i[12], n129);
  or U187 ( n129, n130, add1_i[12]);
  nand U188 ( n120, n122, n123);
  nand U189 ( n122, add1_i[13], n125);
  nand U190 ( n123, add2_i[13], n124);
  or U191 ( n124, n125, add1_i[13]);
  nand U192 ( n115, n117, n118);
  nand U193 ( n117, add1_i[14], n120);
  nand U194 ( n118, add2_i[14], n119);
  or U195 ( n119, n120, add1_i[14]);
  nand U196 ( n110, n112, n113);
  nand U197 ( n112, add1_i[15], n115);
  nand U198 ( n113, add2_i[15], n114);
  or U199 ( n114, n115, add1_i[15]);
  nand U200 ( n105, n107, n108);
  nand U201 ( n107, add1_i[16], n110);
  nand U202 ( n108, add2_i[16], n109);
  or U203 ( n109, n110, add1_i[16]);
  nand U204 ( n100, n102, n103);
  nand U205 ( n102, add1_i[17], n105);
  nand U206 ( n103, add2_i[17], n104);
  or U207 ( n104, n105, add1_i[17]);
  nand U208 ( n95, n97, n98);
  nand U209 ( n97, add1_i[18], n100);
  nand U210 ( n98, add2_i[18], n99);
  or U211 ( n99, n100, add1_i[18]);
  nand U212 ( n90, n92, n93);
  nand U213 ( n92, add1_i[19], n95);
  nand U214 ( n93, add2_i[19], n94);
  or U215 ( n94, n95, add1_i[19]);
  nand U216 ( n85, n87, n88);
  nand U217 ( n87, add1_i[20], n90);
  nand U218 ( n88, add2_i[20], n89);
  or U219 ( n89, n90, add1_i[20]);
  nand U220 ( n80, n82, n83);
  nand U221 ( n82, add1_i[21], n85);
  nand U222 ( n83, add2_i[21], n84);
  or U223 ( n84, n85, add1_i[21]);
  nand U224 ( n75, n77, n78);
  nand U225 ( n77, add1_i[22], n80);
  nand U226 ( n78, add2_i[22], n79);
  or U227 ( n79, n80, add1_i[22]);
  nand U228 ( n70, n72, n73);
  nand U229 ( n72, add1_i[23], n75);
  nand U230 ( n73, add2_i[23], n74);
  or U231 ( n74, n75, add1_i[23]);
  nand U232 ( n65, n67, n68);
  nand U233 ( n67, add1_i[24], n70);
  nand U234 ( n68, add2_i[24], n69);
  or U235 ( n69, n70, add1_i[24]);
  nand U236 ( n60, n62, n63);
  nand U237 ( n62, add1_i[25], n65);
  nand U238 ( n63, add2_i[25], n64);
  or U239 ( n64, n65, add1_i[25]);
  nand U240 ( n55, n57, n58);
  nand U241 ( n57, add1_i[26], n60);
  nand U242 ( n58, add2_i[26], n59);
  or U243 ( n59, n60, add1_i[26]);
  nand U244 ( n50, n52, n53);
  nand U245 ( n52, add1_i[27], n55);
  nand U246 ( n53, add2_i[27], n54);
  or U247 ( n54, n55, add1_i[27]);
  nand U248 ( n45, n47, n48);
  nand U249 ( n47, add1_i[28], n50);
  nand U250 ( n48, add2_i[28], n49);
  or U251 ( n49, n50, add1_i[28]);
  nand U252 ( n40, n42, n43);
  nand U253 ( n42, add1_i[29], n45);
  nand U254 ( n43, add2_i[29], n44);
  or U255 ( n44, n45, add1_i[29]);
  nand U256 ( n35, n37, n38);
  nand U257 ( n37, add1_i[30], n40);
  nand U258 ( n38, add2_i[30], n39);
  or U259 ( n39, n40, add1_i[30]);
  nand U260 ( result_o[32], n32, n33);
  nand U261 ( n32, add1_i[31], n35);
  nand U262 ( n33, add2_i[31], n34);
  or U263 ( n34, n35, add1_i[31]);
  nor U264 ( n30, n26, n27);
  not U265 ( n26, add1_i[7]);
  not U266 ( n27, add2_i[7]);
  or U267 ( result_o[0], add1_i[0], add2_i[0]);
  or U268 ( result_o[1], add1_i[1], add2_i[1]);
  or U269 ( result_o[2], add1_i[2], add2_i[2]);
  or U270 ( result_o[3], add1_i[3], add2_i[3]);
  or U271 ( result_o[4], add1_i[4], add2_i[4]);
  or U272 ( result_o[5], add1_i[5], add2_i[5]);
  or U273 ( result_o[6], add1_i[6], add2_i[6]);
endmodule
