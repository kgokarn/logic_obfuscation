// Verilog File 
module broken_array_multiplier8_aor_enc128.bench (op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,product_o[0],product_o[1],product_o[2],product_o[3],product_o[4],
product_o[5],product_o[6],product_o[7],product_o[8],product_o[9],product_o[10],product_o[11],product_o[12],product_o[13],product_o[14],
product_o[15]);

input op1_i[0],op1_i[1],op1_i[2],op1_i[3],op1_i[4],op1_i[5],op1_i[6],op1_i[7],op2_i[0],
op2_i[1],op2_i[2],op2_i[3],op2_i[4],op2_i[5],op2_i[6],op2_i[7],keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127;


output product_o[0], product_o[1], product_o[2], product_o[3], product_o[4], product_o[5], product_o[6], product_o[7], product_o[8], 
product_o[9], product_o[10], product_o[11], product_o[12], product_o[13], product_o[14], product_o[15];

wire xenc98, xenc112, xenc118, xenc58, n206, n203, xenc7, n223, xenc28, 
n238, n237, xenc0, n230, xenc71, xenc76, n231, n239, n236, n234, 
n258, n257, n256, n254, xenc11, n283, xenc25, xenc52, n279, xenc31, 
n298, n275, n325, n326, n208, n327, n328, xenc67, n348, n330, 
n349, xenc62, n347, n355, n356, n319, xenc94, n312, n296, xenc41, 
n361, n307, n313, n310, n359, xenc73, n384, n385, n386, n383, 
n390, n391, n352, n392, n393, xenc53, n399, n341, xenc125, n373, 
xenc4, n370, n402, n441, n442, n443, xenc35, xenc88, n445, n398, 
n406, xenc16, xenc105, xenc44, n429, xenc91, n468, n465, n417, xenc59, 
n409, n224, n225, n219, n221, n357, n358, xenc50, n401, n463, 
n464, n462, n297, xenc12, n265, n276, n273, xenc48, n333, n289, 
xenc110, xenc99, n466, n455, xenc115, n436, xenc95, xenc114, xenc101, xenc86, 
xenc116, n251, n259, xenc47, xenc18, n282, n262, xenc68, n290, n334, 
xenc32, n295, xenc42, xenc123, n321, xenc78, n335, n336, n291, n292, 
n264, n294, xenc84, n261, n260, xenc9, n263, xenc56, n420, n372, 
n419, xenc63, n421, xenc27, n285, n281, n288, n284, xenc49, xenc64, 
n287, n277, n278, n280, xenc70, n253, n252, n255, xenc106, n375, 
n374, xenc54, n376, xenc46, xenc124, n444, n430, n449, xenc5, xenc108, 
n450, n451, n377, n378, xenc55, n343, n379, n246, n247, n249, 
xenc87, xenc38, n232, n235, n233, n452, xenc83, n437, n438, n454, 
n453, xenc21, n423, n422, xenc2, n424, n473, xenc14, n475, n474, 
n476, n477, xenc39, n478, xenc22, xenc96, n308, xenc102, n309, n311, 
xenc117, xenc74, n408, n446, n448, n447, xenc36, n299, xenc60, xenc122, 
n415, n418, n469, n244, n266, n250, n242, n245, n351, n214, 
n353, xenc10, n329, xenc40, n212, xenc57, n332, n394, xenc61, n216, 
n396, n397, xenc93, n395, n435, xenc65, n403, n364, xenc92, xenc26, 
n204, n318, n340, n428, n360, n306, xenc34, n316, n315, xenc1, 
n317, xenc33, n405, n366, n404, xenc109, n407, n380, xenc29, n342, 
xenc89, n381, n382, xenc8, xenc15, n320, n337, xenc45, n338, n339, 
n368, xenc120, n371, n369, xenc23, xenc37, n271, xenc80, n272, n274, 
n387, xenc127, xenc20, n388, n389, xenc24, n345, n344, xenc119, n346, 
n322, n323, n205, xenc111, xenc100, xenc72, n324, n300, n270, xenc97, 
n433, n432, xenc85, n434, xenc75, n268, n470, n471, xenc30, n472, 
xenc121, xenc13, n314, xenc79, n241, n229, n240, xenc126, n243, n226, 
n227, n228, n425, xenc17, n427, n426, n362, n363, n301, n365, 
n413, n414, n412, n416, n303, n304, n269, xenc69, n305, n207, 
xenc81, xenc3, n222, n460, n457, n481, n482, n479, n480, n456, 
xenc107, n220, xenc43, n486, n485, xenc113, n440, n459, xenc103, xenc104, 
n461, n483, n484, xenc90, n218, n439, n209, n354, xenc66, n302, 
n410, n367, n202, n411, n458, n431, n350, n400, n331, n467, 
n267, n210, n293, n286, n248, xenc6, n213, xenc82, n211, n215, 
xenc77, n487, xenc51, xenc19;

xor g0(xenc118, xenc98, xenc112);
xor g1(n203, xenc58, n206);
xor g2(xenc28, xenc7, n223);
xor g3(xenc0, n238, n237);
xor g4(n237, n230, xenc71);
xor g5(n239, xenc76, n231);
xor g6(n238, n236, n234);
xor g7(product_o[12], n258, n257);
xor g8(n258, n256, n254);
xor g9(xenc25, xenc11, n283);
xor g10(n283, xenc52, n279);
xor g11(n275, xenc31, n298);
xor g12(n208, n325, n326);
xor g13(n325, n327, n328);
xor g14(n330, xenc67, n348);
xor g15(n347, n349, xenc62);
xor g16(n319, n355, n356);
xor g17(n296, xenc94, n312);
xor g18(n307, xenc41, n361);
xor g19(n359, n313, n310);
xor g20(n348, xenc73, n384);
xor g21(n383, n385, n386);
xor g22(n352, n390, n391);
xor g23(n390, n392, n393);
xor g24(n341, xenc53, n399);
xor g25(n355, xenc125, n373);
xor g26(n402, xenc4, n370);
xor g27(n384, n441, n442);
xor g28(n442, n443, xenc35);
xor g29(n398, xenc88, n445);
xor g30(n445, n406, xenc16);
xor g31(n429, xenc105, xenc44);
xor g32(n465, xenc91, n468);
xor g33(n409, n417, xenc59);
nand g34(n219, n224, n225);
or g35(n221, n225, n224);
xnor g36(n356, n357, n358);
xnor g37(n399, xenc50, n401);
xnor g38(n462, n463, n464);
xnor g39(n265, n297, xenc12);
xnor g40(n297, n276, n273);
xnor g41(n289, xenc48, n333);
xnor g42(n333, xenc110, xenc99);
xnor g43(n441, n465, n466);
xnor g44(n436, n455, xenc115);
xnor g45(n455, xenc95, xenc114);
xnor g46(n257, xenc101, xenc86);
xnor g47(n259, xenc116, n251);
xnor g48(n282, xenc47, xenc18);
xnor g49(n290, n262, xenc68);
nand g50(n295, n334, xenc32);
or g51(n334, xenc42, xenc123);
nand g52(n335, n321, xenc78);
nand g53(n336, xenc123, xenc42);
nand g54(n264, n291, n292);
nand g55(n291, xenc48, xenc99);
nand g56(n292, xenc110, n294);
or g57(n294, xenc99, xenc48);
nand g58(n251, xenc84, n261);
nand g59(n260, xenc47, xenc68);
nand g60(n261, n262, xenc9);
or g61(n263, xenc68, xenc47);
nand g62(n372, xenc56, n420);
nand g63(n419, xenc53, n401);
nand g64(n420, xenc50, xenc63);
or g65(n421, n401, xenc53);
nand g66(n281, xenc27, n285);
nand g67(n284, n289, n288);
nand g68(n285, xenc49, xenc64);
or g69(n287, n288, n289);
nand g70(n256, n277, n278);
nand g71(n277, xenc11, xenc52);
nand g72(n278, n279, n280);
or g73(n280, xenc52, xenc11);
nand g74(n236, xenc70, n253);
nand g75(n252, n257, n256);
nand g76(n253, n254, n255);
or g77(n255, n256, n257);
nand g78(n313, xenc106, n375);
nand g79(n374, n355, n358);
nand g80(n375, n357, xenc54);
or g81(n376, n355, n358);
and g82(n444, xenc46, xenc124);
or g83(n449, n429, n430);
nand g84(n450, xenc5, xenc108);
nand g85(n451, n430, n429);
nand g86(n358, n377, n378);
or g87(n377, n341, xenc55);
nand g88(n378, n343, n379);
nand g89(n379, xenc55, n341);
and g90(n230, n246, n247);
nand g91(n246, xenc101, n251);
nand g92(n247, xenc116, n249);
or g93(n249, xenc101, n251);
nand g94(n225, xenc87, xenc38);
nand g95(n232, n237, n236);
nand g96(n233, n234, n235);
or g97(n235, n236, n237);
and g98(n430, n452, xenc83);
or g99(n452, n437, n438);
nand g100(n453, n436, n454);
nand g101(n454, n437, n438);
nand g102(n401, xenc21, n423);
nand g103(n422, n384, n385);
nand g104(n423, n386, xenc2);
or g105(n424, n385, n384);
nand g106(n468, n473, xenc14);
nand g107(n473, xenc105, n464);
nand g108(n474, n463, n475);
or g109(n475, n464, xenc105);
nand g110(n464, n476, n477);
nand g111(n476, xenc95, xenc115);
nand g112(n477, xenc114, xenc39);
or g113(n478, xenc115, xenc95);
and g114(n276, xenc22, xenc96);
nand g115(n308, n312, n313);
nand g116(n309, n310, xenc102);
or g117(n311, n312, n313);
and g118(n408, xenc117, xenc74);
or g119(n446, n441, xenc35);
nand g120(n447, n443, n448);
nand g121(n448, xenc35, n441);
xnor g122(n361, xenc36, n299);
xnor g123(n298, xenc60, xenc122);
xnor g124(n469, n415, n418);
xnor g125(n250, n244, n266);
xnor g126(n266, n242, n245);
xnor g127(n214, n351, n352);
xnor g128(n351, n353, xenc10);
xnor g129(n212, n329, xenc40);
xnor g130(n329, xenc57, n332);
xnor g131(n216, n394, xenc61);
xnor g132(n394, n396, n397);
xnor g133(n395, xenc93, n436);
xnor g134(n435, n437, n438);
xnor g135(n373, xenc65, n403);
xnor g136(n403, n364, xenc92);
xnor g137(n204, xenc26, xenc42);
xnor g138(n318, xenc123, n321);
xnor g139(n326, n340, n341);
xnor g140(n340, xenc55, n343);
xnor g141(n391, n428, n429);
xnor g142(n428, n430, xenc5);
xnor g143(n312, n360, n307);
xnor g144(n360, n306, xenc60);
nand g145(n288, xenc34, n316);
nand g146(n315, n206, xenc58);
nand g147(n316, xenc112, xenc1);
or g148(n317, xenc58, n206);
nand g149(n366, xenc33, n405);
or g150(n404, xenc88, xenc16);
nand g151(n405, n406, xenc109);
nand g152(n407, xenc16, xenc88);
and g153(n342, n380, xenc29);
nand g154(n380, xenc62, n349);
nand g155(n381, n348, xenc89);
or g156(n382, n349, xenc62);
and g157(n320, xenc8, xenc15);
nand g158(n337, n328, n327);
nand g159(n338, n326, xenc45);
or g160(n339, n327, n328);
and g161(n306, n368, xenc120);
nand g162(n368, n373, xenc4);
nand g163(n369, n370, n371);
or g164(n371, xenc4, n373);
and g165(n244, xenc23, xenc37);
or g166(n271, xenc12, n276);
nand g167(n272, n273, xenc80);
nand g168(n274, xenc12, n276);
nand g169(n349, n387, xenc127);
or g170(n387, n353, xenc10);
nand g171(n388, n352, xenc20);
nand g172(n389, n353, xenc10);
nand g173(n327, xenc24, n345);
nand g174(n344, xenc57, n332);
nand g175(n345, xenc40, xenc119);
or g176(n346, xenc57, n332);
nand g177(n205, n322, n323);
or g178(n322, xenc111, xenc100);
nand g179(n323, xenc72, n324);
nand g180(n324, xenc111, xenc100);
nand g181(n270, n299, n300);
nand g182(n300, xenc41, xenc36);
nand g183(n392, xenc97, n433);
or g184(n432, n396, n397);
nand g185(n433, xenc61, xenc85);
nand g186(n434, n396, n397);
and g187(n242, xenc60, xenc75);
nand g188(n268, xenc31, xenc122);
and g189(n417, n470, n471);
nand g190(n470, n466, n468);
nand g191(n471, xenc91, xenc30);
or g192(n472, n468, n466);
xnor g193(xenc13, n289, xenc121);
xnor g194(n314, xenc49, n288);
nand g195(n229, xenc79, n241);
or g196(n240, n245, n244);
nand g197(n241, n242, xenc126);
nand g198(n243, n244, n245);
nand g199(n224, n226, n227);
or g200(n226, n231, n230);
nand g201(n227, n228, xenc76);
nand g202(n228, n230, n231);
nand g203(n385, n425, xenc17);
nand g204(n425, n393, n392);
nand g205(n426, n391, n427);
or g206(n427, n392, n393);
and g207(n301, n362, n363);
nand g208(n362, xenc65, xenc92);
nand g209(n363, n364, n365);
or g210(n365, xenc92, xenc65);
nand g211(n412, n413, n414);
or g212(n413, n418, n417);
nand g213(n414, n415, n416);
nand g214(n416, n417, n418);
and g215(n269, n303, n304);
or g216(n303, n307, n306);
nand g217(n304, xenc60, xenc69);
nand g218(n305, n306, n307);
xnor g219(product_o[8], n207, xenc72);
xnor g220(n207, xenc111, xenc100);
nand g221(n223, op2_i[7], op1_i[7]);
nand g222(n222, xenc81, xenc3);
and g223(n457, op2_i[2], n460, op1_i[2]);
xnor g224(n460, n481, n482);
nand g225(n481, op1_i[3], op2_i[1]);
and g226(n482, op1_i[4], op2_i[0]);
xnor g227(n456, n479, n480);
nand g228(n479, op1_i[4], op2_i[1]);
and g229(n480, op1_i[5], op2_i[0]);
nand g230(product_o[15], xenc3, xenc107);
nand g231(n220, op1_i[7], xenc81, op2_i[7]);
xnor g232(n466, xenc43, n486);
nand g233(n485, op1_i[6], op2_i[1]);
and g234(n486, op1_i[7], op2_i[0]);
xnor g235(n440, xenc113, n460);
nand g236(n459, op1_i[2], op2_i[2]);
xnor g237(n461, xenc103, xenc104);
nand g238(n483, op1_i[5], op2_i[1]);
and g239(n484, op1_i[6], op2_i[0]);
xnor g240(n218, xenc90, n440);
nand g241(n439, op1_i[1], op2_i[3]);
nand g242(n209, op1_i[0], n212, op2_i[7]);
nand g243(n353, op1_i[0], n216, op2_i[5]);
nand g244(n437, op2_i[3], n440, op1_i[1]);
nand g245(n396, op2_i[4], n218, op1_i[0]);
nand g246(n418, op2_i[2], op1_i[6]);
nand g247(n438, op2_i[3], op1_i[2]);
nand g248(n397, op2_i[4], op1_i[1]);
nand g249(n354, op2_i[5], op1_i[1]);
nand g250(n302, op1_i[7], xenc66);
and g251(n367, xenc36, n410);
nand g252(n410, n202, n411);
nand g253(n411, op2_i[2], op1_i[7]);
not g254(n202, xenc66);
and g255(n458, op1_i[3], op2_i[2]);
and g256(n431, op2_i[3], op1_i[3]);
and g257(n393, op2_i[4], op1_i[2]);
and g258(n350, op2_i[5], op1_i[2]);
and g259(n463, op1_i[4], op2_i[2]);
and g260(n415, op2_i[1], op1_i[7]);
and g261(n400, op2_i[4], op1_i[4]);
and g262(n364, op2_i[3], op1_i[6]);
and g263(n331, op2_i[6], op1_i[0], n214);
and g264(n386, op2_i[4], op1_i[3]);
and g265(n467, op1_i[5], op2_i[2]);
and g266(n443, op2_i[3], op1_i[4]);
and g267(n406, op2_i[3], op1_i[5]);
and g268(n267, op2_i[4], op1_i[6]);
nand g269(n245, op2_i[5], op1_i[7]);
nand g270(n210, op2_i[7], op1_i[1]);
and g271(n332, op2_i[6], op1_i[1]);
and g272(n343, op2_i[5], op1_i[3]);
and g273(n299, op2_i[3], op1_i[7]);
and g274(n321, op2_i[6], op1_i[3]);
and g275(n273, op2_i[5], op1_i[6]);
and g276(n328, op2_i[6], op1_i[2]);
and g277(n206, op2_i[7], op1_i[2]);
and g278(n357, op2_i[5], op1_i[4]);
and g279(n293, op2_i[6], op1_i[4]);
and g280(n286, op2_i[7], op1_i[3]);
and g281(n262, op2_i[6], op1_i[5]);
and g282(n248, op2_i[6], op1_i[6]);
xnor g283(product_o[6], xenc6, n214);
nand g284(n213, op2_i[6], op1_i[0]);
xnor g285(product_o[7], xenc82, n212);
nand g286(n211, op2_i[7], op1_i[0]);
and g287(n370, op2_i[4], op1_i[5]);
and g288(n310, op2_i[5], op1_i[5]);
xnor g289(product_o[5], n215, n216);
nand g290(n215, op2_i[5], op1_i[0]);
nand g291(n231, op2_i[6], op1_i[7]);
xnor g292(product_o[4], xenc77, n218);
nand g293(n487, op2_i[4], op1_i[0]);
and g294(n279, op2_i[7], op1_i[4]);
and g295(n254, op2_i[7], op1_i[5]);
and g296(n234, op2_i[7], op1_i[6]);
and g297(xenc51, op2_i[0], op1_i[0]);
and g298(product_o[1], op2_i[1], op1_i[0]);
and g299(xenc19, op2_i[2], op1_i[0]);
and g300(product_o[3], op2_i[3], op1_i[0]);
or g301(product_o[13], xenc0, keyinput0);
or g302(xenc1, n317, keyinput1);
or g303(xenc2, n424, keyinput2);
or g304(xenc3, n219, keyinput3);
or g305(xenc4, n372, keyinput4);
or g306(xenc5, n431, keyinput5);
or g307(xenc6, n213, keyinput6);
or g308(xenc7, n222, keyinput7);
and g309(xenc8, n337, keyinput8);
and g310(xenc9, n263, keyinput9);
or g311(xenc10, n354, keyinput10);
or g312(xenc11, n282, keyinput11);
or g313(xenc12, n275, keyinput12);
or g314(product_o[10], xenc13, keyinput13);
and g315(xenc14, n474, keyinput14);
and g316(xenc15, n338, keyinput15);
and g317(xenc16, n408, keyinput16);
or g318(xenc17, n426, keyinput17);
and g319(xenc18, n290, keyinput18);
or g320(product_o[2], xenc19, keyinput19);
and g321(xenc20, n389, keyinput20);
and g322(xenc21, n422, keyinput21);
or g323(xenc22, n308, keyinput22);
or g324(xenc23, n271, keyinput23);
and g325(xenc24, n344, keyinput24);
or g326(product_o[11], xenc25, keyinput25);
and g327(xenc26, n318, keyinput26);
and g328(xenc27, n284, keyinput27);
or g329(product_o[14], xenc28, keyinput28);
and g330(xenc29, n381, keyinput29);
or g331(xenc30, n472, keyinput30);
and g332(xenc31, n269, keyinput31);
and g333(xenc32, n335, keyinput32);
and g334(xenc33, n404, keyinput33);
or g335(xenc34, n315, keyinput34);
or g336(xenc35, n444, keyinput35);
or g337(xenc36, n302, keyinput36);
and g338(xenc37, n272, keyinput37);
and g339(xenc38, n233, keyinput38);
or g340(xenc39, n478, keyinput39);
and g341(xenc40, n330, keyinput40);
or g342(xenc41, n301, keyinput41);
and g343(xenc42, n319, keyinput42);
and g344(xenc43, n485, keyinput43);
and g345(xenc44, n462, keyinput44);
and g346(xenc45, n339, keyinput45);
and g347(xenc46, n449, keyinput46);
and g348(xenc47, n265, keyinput47);
and g349(xenc48, n296, keyinput48);
and g350(xenc49, n286, keyinput49);
or g351(xenc50, n400, keyinput50);
and g352(product_o[0], xenc51, keyinput51);
and g353(xenc52, n281, keyinput52);
and g354(xenc53, n398, keyinput53);
or g355(xenc54, n376, keyinput54);
and g356(xenc55, n342, keyinput55);
and g357(xenc56, n419, keyinput56);
or g358(xenc57, n331, keyinput57);
and g359(xenc58, n205, keyinput58);
or g360(xenc59, n469, keyinput59);
and g361(xenc60, n267, keyinput60);
or g362(xenc61, n395, keyinput61);
or g363(xenc62, n350, keyinput62);
and g364(xenc63, n421, keyinput63);
or g365(xenc64, n287, keyinput64);
or g366(xenc65, n367, keyinput65);
or g367(xenc66, n412, keyinput66);
and g368(xenc67, n347, keyinput67);
or g369(xenc68, n264, keyinput68);
or g370(xenc69, n305, keyinput69);
or g371(xenc70, n252, keyinput70);
and g372(xenc71, n239, keyinput71);
and g373(xenc72, n208, keyinput72);
and g374(xenc73, n383, keyinput73);
and g375(xenc74, n447, keyinput74);
and g376(xenc75, n268, keyinput75);
and g377(xenc76, n229, keyinput76);
and g378(xenc77, n487, keyinput77);
and g379(xenc78, n336, keyinput78);
and g380(xenc79, n240, keyinput79);
and g381(xenc80, n274, keyinput80);
and g382(xenc81, n221, keyinput81);
and g383(xenc82, n211, keyinput82);
or g384(xenc83, n453, keyinput83);
and g385(xenc84, n260, keyinput84);
and g386(xenc85, n434, keyinput85);
or g387(xenc86, n259, keyinput86);
and g388(xenc87, n232, keyinput87);
or g389(xenc88, n409, keyinput88);
and g390(xenc89, n382, keyinput89);
or g391(xenc90, n439, keyinput90);
or g392(xenc91, n467, keyinput91);
or g393(xenc92, n366, keyinput92);
or g394(xenc93, n435, keyinput93);
or g395(xenc94, n359, keyinput94);
or g396(xenc95, n457, keyinput95);
and g397(xenc96, n309, keyinput96);
and g398(xenc97, n432, keyinput97);
or g399(xenc98, n203, keyinput98);
or g400(xenc99, n295, keyinput99);
or g401(xenc100, n210, keyinput100);
or g402(xenc101, n250, keyinput101);
or g403(xenc102, n311, keyinput102);
or g404(xenc103, n483, keyinput103);
or g405(xenc104, n484, keyinput104);
or g406(xenc105, n461, keyinput105);
or g407(xenc106, n374, keyinput106);
or g408(xenc107, n220, keyinput107);
or g409(xenc108, n451, keyinput108);
and g410(xenc109, n407, keyinput109);
and g411(xenc110, n293, keyinput110);
and g412(xenc111, n209, keyinput111);
and g413(xenc112, n204, keyinput112);
and g414(xenc113, n459, keyinput113);
or g415(xenc114, n458, keyinput114);
and g416(xenc115, n456, keyinput115);
and g417(xenc116, n248, keyinput116);
and g418(xenc117, n446, keyinput117);
or g419(product_o[9], xenc118, keyinput118);
and g420(xenc119, n346, keyinput119);
and g421(xenc120, n369, keyinput120);
and g422(xenc121, n314, keyinput121);
or g423(xenc122, n270, keyinput122);
and g424(xenc123, n320, keyinput123);
or g425(xenc124, n450, keyinput124);
or g426(xenc125, n402, keyinput125);
or g427(xenc126, n243, keyinput126);
or g428(xenc127, n388, keyinput127);
endmodule
