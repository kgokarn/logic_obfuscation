module xnor_based_ripple_carry_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110;

  xor U56 ( result_o[9], add2_i[9], n51);
  xor U57 ( result_o[8], add2_i[8], n52);
  xor U58 ( result_o[7], add2_i[7], n53);
  xor U59 ( result_o[6], add2_i[6], n54);
  xor U60 ( result_o[5], n55, add2_i[5]);
  xor U61 ( result_o[4], n56, add2_i[4]);
  xor U62 ( result_o[15], add2_i[15], n65);
  xor U63 ( n65, n66, add1_i[15]);
  xor U64 ( result_o[14], add2_i[14], n69);
  xor U65 ( n69, n70, add1_i[14]);
  xor U66 ( result_o[13], add2_i[13], n73);
  xor U67 ( n73, n74, add1_i[13]);
  xor U68 ( result_o[12], add2_i[12], n77);
  xor U69 ( n77, n78, add1_i[12]);
  xor U70 ( result_o[11], add2_i[11], n81);
  xor U71 ( n81, n82, add1_i[11]);
  xor U72 ( result_o[10], add2_i[10], n85);
  xor U73 ( n85, n86, add1_i[10]);
  xor U74 ( n51, n89, add1_i[9]);
  xor U75 ( n52, n92, add1_i[8]);
  xor U76 ( n53, n95, add1_i[7]);
  xor U77 ( n54, n98, add1_i[6]);
  xor U78 ( n55, n101, add1_i[5]);
  xor U79 ( n56, n104, add1_i[4]);
  xor U80 ( n62, add1_i[1], add2_i[1]);
  xor U81 ( n59, add1_i[2], add2_i[2]);
  xor U82 ( n57, add1_i[3], add2_i[3]);
  nor U83 ( result_o[1], n61, n62);
  nor U84 ( result_o[3], n47, n57);
  not U85 ( n47, n58);
  nor U86 ( result_o[2], n48, n59);
  not U87 ( n48, n60);
  nor U88 ( n61, n50, add1_i[0]);
  not U89 ( n50, result_o[0]);
  xnor U90 ( result_o[0], add1_i[0], add2_i[0]);
  nand U91 ( n104, n105, n106);
  nand U92 ( n105, add1_i[3], add2_i[3]);
  nand U93 ( n106, n57, n58);
  nand U94 ( n60, n109, n110);
  nand U95 ( n109, add1_i[1], add2_i[1]);
  nand U96 ( n110, n62, n49);
  not U97 ( n49, n61);
  nand U98 ( n58, n107, n108);
  nand U99 ( n107, add1_i[2], add2_i[2]);
  nand U100 ( n108, n59, n60);
  nand U101 ( n82, n83, n84);
  nand U102 ( n83, add1_i[10], n86);
  nand U103 ( n84, add2_i[10], n85);
  nand U104 ( n78, n79, n80);
  nand U105 ( n79, add1_i[11], n82);
  nand U106 ( n80, add2_i[11], n81);
  nand U107 ( n74, n75, n76);
  nand U108 ( n75, add1_i[12], n78);
  nand U109 ( n76, add2_i[12], n77);
  nand U110 ( n70, n71, n72);
  nand U111 ( n71, add1_i[13], n74);
  nand U112 ( n72, add2_i[13], n73);
  nand U113 ( n66, n67, n68);
  nand U114 ( n67, add1_i[14], n70);
  nand U115 ( n68, add2_i[14], n69);
  nand U116 ( n98, n99, n100);
  nand U117 ( n99, add1_i[5], n101);
  nand U118 ( n100, add2_i[5], n55);
  nand U119 ( n95, n96, n97);
  nand U120 ( n96, add1_i[6], n98);
  nand U121 ( n97, add2_i[6], n54);
  nand U122 ( n92, n93, n94);
  nand U123 ( n93, add1_i[7], n95);
  nand U124 ( n94, add2_i[7], n53);
  nand U125 ( n89, n90, n91);
  nand U126 ( n90, add1_i[8], n92);
  nand U127 ( n91, add2_i[8], n52);
  nand U128 ( n86, n87, n88);
  nand U129 ( n87, add1_i[9], n89);
  nand U130 ( n88, add2_i[9], n51);
  nand U131 ( n101, n102, n103);
  nand U132 ( n102, add1_i[4], n104);
  nand U133 ( n103, add2_i[4], n56);
  nand U134 ( result_o[16], n63, n64);
  nand U135 ( n63, add1_i[15], n66);
  nand U136 ( n64, add2_i[15], n65);
endmodule
