// Verilog File 
module xnor_based_ripple_carry_adder32_aor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire xenc23, xenc72, n203, n331, xenc76, n228, xenc119, n237, xenc58, 
xenc40, n250, xenc33, xenc96, xenc92, xenc86, n288, xenc116, n292, xenc113, 
n296, xenc71, n190, n199, n216, n267, xenc42, xenc98, n326, xenc105, 
n327, n328, n217, xenc35, n218, n325, n329, n340, n274, xenc101, 
xenc77, n201, n322, xenc14, n339, n179, xenc57, xenc6, xenc109, n313, 
xenc66, xenc12, n335, xenc16, n320, xenc2, xenc90, n249, xenc79, xenc110, 
xenc43, xenc107, xenc74, xenc61, xenc25, xenc9, n255, n233, xenc87, xenc18, 
xenc121, xenc83, n343, n342, n346, xenc13, n330, n332, xenc7, xenc95, 
n333, n268, n334, xenc31, xenc48, n270, xenc111, n336, n212, xenc50, 
n337, xenc85, xenc102, n338, n269, xenc103, n232, n341, n264, xenc49, 
n263, n242, n241, xenc19, n344, xenc84, n345, n238, n350, xenc60, 
xenc126, n347, n349, n348, n276, n285, xenc82, n284, xenc15, xenc97, 
n351, n352, xenc22, xenc123, n281, n280, n367, n353, n362, n355, 
n354, n356, xenc41, xenc118, n260, n297, xenc106, xenc46, n210, n357, 
n361, n358, n360, n234, xenc36, n359, xenc29, xenc65, n206, xenc100, 
n215, xenc55, n214, xenc67, n183, n193, n181, n189, xenc54, xenc38, 
n191, xenc69, xenc17, xenc59, n366, n365, n195, n200, n319, n222, 
n178, n221, xenc4, xenc117, xenc20, n363, n315, n321, n364, xenc80, 
xenc24, n272, n186, xenc10, xenc62, n196, n198, n265, xenc127, xenc45, 
n266, n305, xenc39, n304, n239, xenc108, xenc51, n309, xenc112, xenc52, 
n187, xenc89, n301, n300, n316, n312, xenc21, n318, n317, n324, 
n323, n368, n202, n369, xenc63, xenc0, xenc68, n290, n298, n307, 
xenc37, xenc32, xenc3, n220, xenc122, n294, n293, xenc115, n303, n244, 
n243, n245, n261, xenc73, n231, n246, n275, n273, xenc81, n204, 
xenc114, n208, n253, n279, n278, n277, n207, n211, xenc64, xenc47, 
n256, n283, xenc28, n282, n306, n302, n314, n188, n235, xenc94, 
n248, n251, n286, xenc70, xenc5, xenc104, n311, xenc30, xenc88, xenc44, 
n180, n219, xenc34, n229, n226, xenc91, xenc8, n252, xenc93, n291, 
xenc75, n289, xenc56, n192, xenc99, xenc27, xenc1, n205, n197, xenc53, 
n225, n227, n223, xenc26, n224, n258, n257, xenc78, xenc124, n259, 
n299, xenc11, n310, xenc125, n209, n213, n230, n236, xenc120, n240, 
n254, n262, n287, n295, n308;

xor g0(xenc72, add2_i[8], xenc23);
xor g1(n203, add2_i[3], add1_i[3]);
xor g2(result_o[29], add2_i[29], n331);
xor g3(xenc119, xenc76, n228);
xor g4(xenc58, n237, add2_i[25]);
xor g5(result_o[24], xenc40, add2_i[24]);
xor g6(xenc33, add2_i[22], n250);
xor g7(result_o[16], add2_i[16], xenc96);
xor g8(xenc86, xenc92, add2_i[15]);
xor g9(xenc116, add2_i[14], n288);
xor g10(xenc113, add2_i[13], n292);
xor g11(result_o[12], add2_i[12], n296);
xor g12(result_o[10], add2_i[10], xenc71);
xor g13(n190, add1_i[7], add2_i[7]);
xor g14(n199, add1_i[4], add2_i[4]);
xor g15(n216, add1_i[2], add2_i[2]);
xor g16(n267, add1_i[0], add2_i[0]);
xnor g17(n326, xenc42, xenc98);
not g18(n327, xenc105);
not g19(n328, n327);
or g20(n325, n217, xenc35, n218);
nand g21(n340, n329, add1_i[18]);
not g22(n329, n274);
nand g23(n322, xenc101, xenc77, n201);
nand g24(n339, xenc14, add2_i[17], add1_i[18]);
nand g25(n313, n179, xenc57, xenc6, xenc109);
and g26(n335, xenc66, add2_i[18], xenc12);
nand g27(n320, xenc16, add2_i[5], add1_i[5]);
nand g28(n249, xenc2, xenc90, add2_i[22]);
xor g29(xenc110, add2_i[9], xenc79);
xor g30(xenc107, add2_i[11], xenc43);
xor g31(xenc74, add2_i[17], xenc14);
xor g32(xenc25, add2_i[19], xenc61);
xor g33(result_o[20], add2_i[20], xenc9);
xor g34(result_o[21], add2_i[21], n255);
xor g35(xenc87, add2_i[26], n233);
xor g36(xenc18, add2_i[30], n328);
xor g37(xenc83, xenc121, add2_i[31]);
not g38(n343, add1_i[24]);
not g39(n342, add1_i[19]);
not g40(n346, add1_i[25]);
not g41(n330, xenc13);
not g42(n331, n330);
and g43(n332, xenc57, xenc6);
nand g44(n333, xenc7, xenc95);
and g45(n268, add1_i[1], add2_i[1]);
or g46(n334, add1_i[0], add2_i[0]);
nand g47(n270, xenc31, xenc48);
or g48(n336, xenc111, add1_i[18]);
nand g49(n337, n212, xenc50);
nand g50(n338, xenc85, xenc102);
and g51(n269, xenc66, xenc12);
nand g52(n341, xenc103, n232);
xnor g53(n263, n264, xenc49);
xnor g54(n241, n242, n343);
not g55(n344, xenc19);
not g56(n345, xenc84);
xnor g57(n237, n238, n346);
not g58(n350, add1_i[13]);
nor g59(n217, xenc60, xenc126);
xor g60(n347, n242, add1_i[24]);
not g61(n349, add1_i[15]);
not g62(n348, add1_i[17]);
xnor g63(n276, xenc42, xenc98);
xnor g64(n284, n285, xenc82);
xnor g65(n292, xenc15, xenc97);
not g66(n351, add1_i[14]);
not g67(n352, add1_i[16]);
xnor g68(n288, xenc22, xenc123);
xnor g69(n280, n281, n352);
nor g70(n353, add1_i[0], add2_i[0], n367);
not g71(n362, add1_i[29]);
not g72(n355, add1_i[12]);
not g73(n354, add1_i[20]);
not g74(n356, add1_i[30]);
xnor g75(n260, xenc41, xenc118);
xnor g76(n296, n297, n355);
xnor g77(n210, xenc106, xenc46);
xor g78(n357, add1_i[6], add2_i[6]);
not g79(n361, add1_i[21]);
not g80(n358, add1_i[26]);
not g81(n360, add1_i[31]);
xnor g82(n233, n234, xenc36);
xnor g83(n359, add1_i[2], add2_i[2]);
xnor g84(n206, xenc29, xenc65);
xnor g85(n255, xenc100, n361);
xnor g86(n214, n215, xenc55);
not g87(n183, xenc67);
not g88(n181, n193);
nor g89(xenc38, n189, xenc54);
nor g90(n189, n191, xenc69);
nor g91(xenc59, xenc77, xenc17, xenc67);
not g92(result_o[0], n267);
not g93(n366, add1_i[11]);
not g94(n365, add1_i[9]);
xor g95(n195, add1_i[6], add2_i[6]);
xnor g96(n193, add1_i[5], add2_i[5]);
nor g97(n218, add2_i[1], add1_i[1]);
nor g98(n200, add2_i[3], add1_i[3]);
nand g99(n319, add1_i[6], add2_i[6]);
nand g100(n221, n222, n178);
xnor g101(n228, add2_i[28], n178);
xor g102(xenc20, xenc4, xenc117);
xor g103(n363, add1_i[23], add2_i[23]);
and g104(n250, xenc90, xenc2);
nand g105(n315, add2_i[7], add1_i[7]);
nand g106(n321, add1_i[4], add2_i[4]);
xnor g107(xenc80, add2_i[18], n364);
nand g108(n364, xenc24, n272);
not g109(n178, add1_i[28]);
not g110(n186, add2_i[27]);
nor g111(n196, xenc10, xenc62);
and g112(n198, add1_i[5], add2_i[5]);
nor g113(xenc45, n265, xenc127);
nor g114(n265, n367, n218);
nor g115(n266, add1_i[0], n267);
and g116(n304, n305, xenc39);
nand g117(n239, add1_i[24], n242);
nand g118(n309, xenc108, xenc51);
xnor g119(n187, xenc112, xenc52);
xnor g120(n300, xenc89, n301);
and g121(n367, add1_i[1], add2_i[1]);
nand g122(n312, xenc109, n316);
not g123(n179, xenc69);
nand g124(n316, xenc54, xenc21);
nand g125(n317, n179, n318);
and g126(n368, n324, n323);
and g127(n369, n202, n323);
nand g128(n324, add1_i[2], add2_i[2]);
nand g129(n323, add2_i[3], add1_i[3]);
and g130(n202, xenc63, n324);
nor g131(xenc68, n202, xenc0);
nand g132(n201, xenc63, n368);
nand g133(n212, add1_i[29], n215);
nand g134(n290, xenc15, add1_i[13]);
nand g135(n298, add1_i[11], n301);
nand g136(n307, xenc112, add1_i[9]);
nand g137(n215, xenc37, xenc32);
nand g138(n220, add2_i[28], xenc3);
nand g139(n293, xenc122, n294);
nand g140(n301, xenc115, xenc39);
nand g141(n303, add2_i[10], xenc71);
nand g142(n242, n244, n243);
nand g143(n244, n245, add2_i[23]);
or g144(n272, xenc111, add1_i[18]);
nand g145(n264, n270, xenc24);
nand g146(n261, add1_i[19], n264);
nand g147(n231, add1_i[26], xenc73);
nand g148(n246, n249, xenc2);
nand g149(n273, n275, n274);
nand g150(n274, add1_i[17], xenc42);
nand g151(n204, add1_i[31], xenc81);
nand g152(n208, add1_i[30], xenc114);
nand g153(n253, add1_i[21], xenc100);
nand g154(n277, n279, n278);
nand g155(n207, xenc7, xenc95);
nand g156(n211, n212, xenc50);
nand g157(n234, xenc85, xenc102);
nand g158(n256, xenc64, xenc47);
nand g159(n281, n283, xenc28);
nand g160(n282, n285, add1_i[15]);
or g161(n305, n306, add1_i[10]);
nand g162(n302, add1_i[10], n306);
xnor g163(n188, n314, add1_i[8]);
nand g164(n235, add1_i[25], n238);
nand g165(n248, add1_i[22], xenc94);
or g166(n251, xenc94, add1_i[22]);
nand g167(n286, add1_i[14], xenc22);
nand g168(n294, add1_i[12], n297);
nand g169(n306, xenc70, xenc5);
nand g170(n311, xenc104, n313, add1_i[8]);
nand g171(n314, n313, xenc104);
nor g172(xenc30, n196, n357);
xnor g173(xenc44, add2_i[27], xenc88);
not g174(n180, n357);
nand g175(n219, add1_i[28], xenc76);
or g176(n229, xenc88, xenc34);
nand g177(n226, xenc103, n232);
nand g178(n238, n239, xenc91);
nand g179(n252, xenc8, n253);
nand g180(n285, xenc93, n286);
nand g181(n289, n291, xenc75);
nand g182(n318, xenc56, n357);
nand g183(n192, n319, n320);
nand g184(result_o[32], xenc99, xenc27);
nor g185(xenc1, n332, xenc56);
nand g186(n205, add2_i[31], xenc121);
nor g187(n197, n332, n193);
nor g188(n191, n193, n332, xenc53);
nand g189(n227, n229, n225);
nand g190(n222, n223, xenc26);
nand g191(n224, n225, xenc34);
nand g192(n243, add1_i[23], xenc117);
or g193(n245, xenc117, add1_i[23]);
nand g194(n258, add1_i[20], xenc41);
nand g195(n257, add2_i[20], xenc9);
nand g196(n259, xenc78, xenc124);
nand g197(n278, add1_i[16], n281);
nand g198(n283, add2_i[15], xenc92);
nand g199(n297, n299, xenc11);
nand g200(n310, xenc19, add2_i[8]);
nor g201(xenc125, n216, n353, n218);
nand g202(n209, add2_i[30], xenc105);
nand g203(n213, add2_i[29], xenc13);
or g204(n223, n341, add1_i[27]);
nand g205(n225, add1_i[27], n341);
xnor g206(n230, n226, add1_i[27]);
nand g207(n232, add2_i[26], n233);
nand g208(n236, add2_i[25], n237);
nand g209(n240, xenc120, add2_i[24]);
nand g210(n254, n255, add2_i[21]);
nand g211(n262, add2_i[19], xenc61);
nand g212(n275, n276, add2_i[17]);
nand g213(n279, xenc96, add2_i[16]);
nand g214(n287, add2_i[14], n288);
nand g215(n291, add2_i[13], n292);
nand g216(n295, add2_i[12], n296);
nand g217(n299, add2_i[11], xenc43);
nand g218(n308, add2_i[9], xenc79);
and g219(xenc0, n203, keyinput0);
and g220(result_o[5], xenc1, keyinput1);
or g221(xenc2, n248, keyinput2);
and g222(xenc3, n221, keyinput3);
and g223(xenc4, n363, keyinput4);
and g224(xenc5, n307, keyinput5);
and g225(xenc6, n322, keyinput6);
and g226(xenc7, n209, keyinput7);
or g227(xenc8, n254, keyinput8);
or g228(xenc9, n260, keyinput9);
or g229(xenc10, n197, keyinput10);
or g230(xenc11, n298, keyinput11);
or g231(xenc12, n340, keyinput12);
and g232(xenc13, n214, keyinput13);
or g233(xenc14, n326, keyinput14);
and g234(xenc15, n293, keyinput15);
or g235(xenc16, n195, keyinput16);
and g236(xenc17, n369, keyinput17);
or g237(result_o[30], xenc18, keyinput18);
and g238(xenc19, n188, keyinput19);
and g239(result_o[23], xenc20, keyinput20);
and g240(xenc21, n317, keyinput21);
and g241(xenc22, n289, keyinput22);
and g242(xenc23, n345, keyinput23);
and g243(xenc24, n269, keyinput24);
and g244(result_o[19], xenc25, keyinput25);
and g245(xenc26, n224, keyinput26);
and g246(xenc27, n205, keyinput27);
or g247(xenc28, n282, keyinput28);
and g248(xenc29, n207, keyinput29);
or g249(result_o[6], xenc30, keyinput30);
and g250(xenc31, n336, keyinput31);
and g251(xenc32, n220, keyinput32);
and g252(result_o[22], xenc33, keyinput33);
and g253(xenc34, n186, keyinput34);
and g254(xenc35, n359, keyinput35);
or g255(xenc36, n358, keyinput36);
and g256(xenc37, n219, keyinput37);
and g257(result_o[7], xenc38, keyinput38);
and g258(xenc39, n302, keyinput39);
and g259(xenc40, n347, keyinput40);
or g260(xenc41, n259, keyinput41);
or g261(xenc42, n277, keyinput42);
or g262(xenc43, n300, keyinput43);
and g263(result_o[27], xenc44, keyinput44);
or g264(result_o[1], xenc45, keyinput45);
or g265(xenc46, n356, keyinput46);
or g266(xenc47, n258, keyinput47);
or g267(xenc48, n335, keyinput48);
and g268(xenc49, n342, keyinput49);
and g269(xenc50, n213, keyinput50);
or g270(xenc51, n311, keyinput51);
or g271(xenc52, n365, keyinput52);
and g272(xenc53, n180, keyinput53);
or g273(xenc54, n190, keyinput54);
or g274(xenc55, n362, keyinput55);
and g275(xenc56, n181, keyinput56);
and g276(xenc57, n321, keyinput57);
and g277(result_o[25], xenc58, keyinput58);
and g278(result_o[4], xenc59, keyinput59);
and g279(xenc60, n334, keyinput60);
or g280(xenc61, n263, keyinput61);
and g281(xenc62, n198, keyinput62);
and g282(xenc63, n325, keyinput63);
and g283(xenc64, n257, keyinput64);
and g284(xenc65, n360, keyinput65);
and g285(xenc66, n339, keyinput66);
or g286(xenc67, n200, keyinput67);
or g287(result_o[3], xenc68, keyinput68);
and g288(xenc69, n192, keyinput69);
or g289(xenc70, n308, keyinput70);
or g290(xenc71, n304, keyinput71);
or g291(result_o[8], xenc72, keyinput72);
or g292(xenc73, n338, keyinput73);
and g293(result_o[17], xenc74, keyinput74);
or g294(xenc75, n290, keyinput75);
and g295(xenc76, n227, keyinput76);
or g296(xenc77, n199, keyinput77);
or g297(xenc78, n261, keyinput78);
or g298(xenc79, n187, keyinput79);
or g299(result_o[18], xenc80, keyinput80);
or g300(xenc81, n333, keyinput81);
or g301(xenc82, n349, keyinput82);
and g302(result_o[31], xenc83, keyinput83);
or g303(xenc84, n344, keyinput84);
and g304(xenc85, n235, keyinput85);
and g305(result_o[15], xenc86, keyinput86);
or g306(result_o[26], xenc87, keyinput87);
and g307(xenc88, n230, keyinput88);
and g308(xenc89, n366, keyinput89);
or g309(xenc90, n251, keyinput90);
and g310(xenc91, n240, keyinput91);
or g311(xenc92, n284, keyinput92);
or g312(xenc93, n287, keyinput93);
and g313(xenc94, n252, keyinput94);
or g314(xenc95, n208, keyinput95);
and g315(xenc96, n280, keyinput96);
and g316(xenc97, n350, keyinput97);
and g317(xenc98, n348, keyinput98);
or g318(xenc99, n204, keyinput99);
and g319(xenc100, n256, keyinput100);
and g320(xenc101, n183, keyinput101);
and g321(xenc102, n236, keyinput102);
and g322(xenc103, n231, keyinput103);
or g323(xenc104, n312, keyinput104);
and g324(xenc105, n210, keyinput105);
or g325(xenc106, n211, keyinput106);
or g326(result_o[11], xenc107, keyinput107);
or g327(xenc108, n310, keyinput108);
and g328(xenc109, n315, keyinput109);
and g329(result_o[9], xenc110, keyinput110);
and g330(xenc111, n273, keyinput111);
or g331(xenc112, n309, keyinput112);
or g332(result_o[13], xenc113, keyinput113);
or g333(xenc114, n337, keyinput114);
and g334(xenc115, n303, keyinput115);
and g335(result_o[14], xenc116, keyinput116);
or g336(xenc117, n246, keyinput117);
and g337(xenc118, n354, keyinput118);
and g338(result_o[28], xenc119, keyinput119);
or g339(xenc120, n241, keyinput120);
or g340(xenc121, n206, keyinput121);
or g341(xenc122, n295, keyinput122);
and g342(xenc123, n351, keyinput123);
or g343(xenc124, n262, keyinput124);
or g344(result_o[2], xenc125, keyinput125);
and g345(xenc126, n268, keyinput126);
or g346(xenc127, n266, keyinput127);
endmodule
