// Verilog File 
module almost_correct_adder32_aor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n262, n263, xenc19, xenc12, xenc100, n269, xenc16, n274, xenc66, 
n287, xenc28, n291, xenc119, n294, n295, n298, xenc102, xenc37, n299, 
xenc40, n317, n302, n321, xenc35, xenc61, n327, xenc53, n339, n351, 
n352, xenc86, xenc43, xenc113, xenc9, n356, n365, n366, n375, xenc62, 
xenc8, n376, n379, n380, xenc127, n389, n390, xenc97, xenc73, n400, 
xenc122, n404, xenc33, xenc13, xenc90, n413, xenc57, n415, xenc27, n424, 
n425, xenc118, xenc104, n429, n436, n437, xenc55, n447, xenc93, n450, 
xenc121, xenc70, n451, xenc51, xenc42, xenc84, n460, xenc39, n472, xenc108, 
n479, n480, xenc109, n485, xenc85, n228, n378, n223, n354, n218, 
n398, xenc126, n402, n410, n394, n409, xenc81, xenc3, n412, n406, 
n411, n374, xenc30, n386, n370, n385, xenc20, n387, xenc47, xenc88, 
n350, n361, n362, n344, xenc44, n363, xenc63, n358, xenc101, n220, 
n340, xenc117, n244, n439, n240, n417, n235, n230, n225, xenc25, 
n243, xenc2, n238, n427, n233, n253, n219, xenc80, n293, n290, 
xenc41, xenc15, n349, n463, n464, n465, n454, xenc74, n466, xenc124, 
n241, n468, n469, n467, xenc6, xenc56, xenc23, xenc59, n442, xenc5, 
xenc94, n443, n445, n440, n444, xenc18, n392, n421, xenc77, n420, 
n384, n422, n423, n418, n395, n368, n396, n359, xenc106, xenc38, 
xenc120, n397, n334, n371, n341, n372, xenc24, n332, xenc68, n369, 
n373, n458, xenc26, n462, n489, xenc49, n491, xenc7, n221, n261, 
xenc83, n259, n234, xenc78, xenc58, xenc31, n229, xenc111, n231, n388, 
n255, xenc48, xenc67, n226, n364, n453, n492, n264, xenc4, xenc45, 
xenc36, n449, n456, n441, n455, xenc0, n457, xenc115, n433, xenc32, 
n432, n434, n431, n266, xenc54, n245, n478, n419, n407, n383, 
n330, xenc79, n320, n318, n475, n476, n474, n477, n278, n279, 
n276, n483, n487, n281, n283, n284, xenc125, n250, n482, n315, 
xenc11, n331, n333, n277, n382, n251, xenc17, n329, n246, n242, 
n488, n249, n288, n272, n247, n237, n232, n227, n222, n267, 
n248, n308, xenc71, n306, xenc64, n310, n309, n325, n342, n289, 
n286, xenc87, xenc82, n337, n345, xenc96, n346, n348, xenc46, n347, 
n296, n297, xenc105, xenc91, n301, n300, xenc98, n252, xenc29, n323, 
n322, n324, xenc103, xenc92, n307, n335, xenc114, n336, xenc21, n313, 
n311, n312, n303, n304, xenc95, xenc76, n305, n490, n282, xenc60, 
n314, n408, n360, n393, xenc75, n484, n486, xenc123, n446, n448, 
n426, n416, n414, xenc10, n401, n399, xenc69, n391, xenc52, xenc72, 
n377, xenc1, n367, n353, n217, n338, n265, xenc34, n459, xenc14, 
n461, n275, n273, n430, n428, xenc65, n405, n403, xenc107, xenc110, 
n381, n357, n355, n328, n326, xenc99, xenc112, n452, xenc50, n481, 
n471, n473, xenc89, n316, n319, n280, n270, n292, n435, n285, 
n343, n239, n236, n224, n470, n260, n257, n258, n256, n254, 
xenc116, n438, xenc22, n268, n271, n493;

xor g0(result_o[9], n262, n263);
xor g1(n263, add2_i[9], add1_i[9]);
xor g2(xenc100, xenc19, xenc12);
xor g3(n269, add2_i[8], add1_i[8]);
xor g4(result_o[7], xenc16, n274);
xor g5(n274, add2_i[7], add1_i[7]);
xor g6(result_o[6], xenc66, n287);
xor g7(n287, add2_i[6], add1_i[6]);
xor g8(xenc119, xenc28, n291);
xor g9(n291, add2_i[5], add1_i[5]);
xor g10(result_o[4], n294, n295);
xor g11(n295, add2_i[4], add1_i[4]);
xor g12(xenc37, n298, xenc102);
xor g13(n299, add2_i[3], add1_i[3]);
xor g14(result_o[30], xenc40, n317);
xor g15(result_o[2], n302, n321);
xor g16(n321, add2_i[2], add1_i[2]);
xor g17(result_o[29], xenc35, xenc61);
xor g18(n327, add2_i[29], add1_i[29]);
xor g19(result_o[28], xenc53, n339);
xor g20(n339, add2_i[28], add1_i[28]);
xor g21(xenc86, n351, n352);
xor g22(n352, add2_i[27], add1_i[27]);
xor g23(xenc9, xenc43, xenc113);
xor g24(n356, add2_i[26], add1_i[26]);
xor g25(result_o[25], n365, n366);
xor g26(n366, add2_i[25], add1_i[25]);
xor g27(xenc8, n375, xenc62);
xor g28(n376, add2_i[24], add1_i[24]);
xor g29(xenc127, n379, n380);
xor g30(n380, add2_i[23], add1_i[23]);
xor g31(result_o[22], n389, n390);
xor g32(n390, add2_i[22], add1_i[22]);
xor g33(result_o[21], xenc97, xenc73);
xor g34(n400, add2_i[21], add1_i[21]);
xor g35(result_o[20], xenc122, n404);
xor g36(n404, add2_i[20], add1_i[20]);
xor g37(xenc90, xenc33, xenc13);
xor g38(n413, add2_i[1], add1_i[1]);
xor g39(xenc27, xenc57, n415);
xor g40(n415, add2_i[19], add1_i[19]);
xor g41(result_o[18], n424, n425);
xor g42(n425, add2_i[18], add1_i[18]);
xor g43(result_o[17], xenc118, xenc104);
xor g44(n429, add2_i[17], add1_i[17]);
xor g45(result_o[16], n436, n437);
xor g46(n437, add2_i[16], add1_i[16]);
xor g47(xenc93, xenc55, n447);
xor g48(n447, add2_i[15], add1_i[15]);
xor g49(xenc70, n450, xenc121);
xor g50(n451, add2_i[14], add1_i[14]);
xor g51(xenc84, xenc51, xenc42);
xor g52(n460, add2_i[13], add1_i[13]);
xor g53(xenc108, xenc39, n472);
xor g54(result_o[11], n479, n480);
xor g55(result_o[10], xenc109, n485);
xor g56(n485, add2_i[10], add1_i[10]);
not g57(n228, xenc85);
not g58(n223, n378);
not g59(n218, n354);
nor g60(n402, n398, xenc126);
and g61(n409, n410, n394);
nand g62(n410, xenc81, xenc3);
nand g63(n411, n412, n406);
nor g64(n378, n374, xenc30);
and g65(n385, n386, n370);
nand g66(n386, xenc20, n387);
nand g67(n387, xenc47, xenc88);
nor g68(n354, n350, n361);
and g69(n361, n362, n344);
nand g70(n362, xenc44, n363);
nand g71(n363, xenc63, n358);
nand g72(n340, xenc101, n220);
not g73(n220, xenc44);
not g74(n244, xenc117);
not g75(n240, n439);
not g76(n235, n417);
not g77(n230, xenc81);
not g78(n225, xenc20);
not g79(n243, xenc25);
not g80(n238, xenc2);
not g81(n233, n427);
nor g82(n350, n253, n219);
nand g83(n290, xenc80, n293);
nand g84(n293, n294, xenc41);
nand g85(n349, n350, xenc15);
nor g86(n454, n463, n464, n465);
nor g87(n439, xenc74, n466);
and g88(n466, xenc124, n241);
nand g89(n467, n468, n469);
or g90(n469, xenc6, n463);
nor g91(n417, n412, xenc56);
and g92(n442, xenc23, xenc59);
nand g93(n443, xenc5, xenc94);
nand g94(n444, n445, n440);
nor g95(n392, xenc47, xenc18);
and g96(n420, n421, xenc77);
nand g97(n421, n384, n422);
nand g98(n422, n423, n418);
nor g99(n368, xenc63, n395);
and g100(n395, n396, n359);
nand g101(n396, xenc106, xenc38);
nand g102(n397, n398, xenc120);
nor g103(n341, n334, n371);
and g104(n371, n372, xenc24);
nand g105(n372, n332, xenc68);
nand g106(n373, n374, n369);
nor g107(n462, n458, xenc26);
nor g108(n491, n489, xenc49);
nor g109(n334, xenc7, n221);
nor g110(n445, n261, xenc83);
nor g111(n423, n259, n234);
nor g112(n412, xenc78, xenc58);
nor g113(n398, xenc31, n229);
nor g114(n388, xenc111, n231);
nor g115(n374, n255, xenc48);
nor g116(n364, xenc67, n226);
nor g117(n264, n453, n492);
nor g118(n492, xenc4, xenc45);
nor g119(n449, n445, xenc36);
and g120(n455, n456, n441);
nand g121(n456, n439, xenc0);
nand g122(n457, n458, n454);
nor g123(n427, n423, xenc115);
and g124(n432, n433, xenc32);
nand g125(n433, n417, n434);
nand g126(n434, xenc74, n431);
nand g127(n478, n266, xenc54, n245);
nand g128(n441, n261, xenc83);
nand g129(n419, n259, n234);
nand g130(n394, xenc31, n229);
nand g131(n370, n255, xenc48);
nand g132(n344, n253, n219);
nand g133(n407, xenc78, xenc58);
nand g134(n383, xenc111, n231);
nand g135(n359, xenc67, n226);
nand g136(n330, xenc7, n221);
nor g137(n318, xenc79, n320);
nor g138(n474, n475, n476);
nor g139(n475, n477, n465, xenc117);
nor g140(n276, n278, n279);
nand g141(n281, n483, n487);
nand g142(n487, n283, n284, xenc125);
not g143(n250, xenc80);
nand g144(n476, xenc6, n482);
or g145(n482, xenc25, n465);
and g146(n320, n315, xenc11);
nand g147(n333, xenc101, n331, n334);
and g148(n277, n283, n284, xenc41);
and g149(n431, n440, xenc59, n441);
and g150(n406, n418, xenc77, xenc32);
and g151(n382, xenc120, n359, n394);
and g152(n358, n369, xenc24, n370);
not g153(n251, n278);
and g154(n329, xenc15, xenc17, n344);
not g155(n245, n489);
not g156(n246, xenc45);
not g157(n242, n468);
not g158(n241, n464);
and g159(n483, n477, n488);
nand g160(n488, n249, n284);
not g161(n249, n288);
not g162(n247, n272);
not g163(n237, xenc5);
not g164(n232, n384);
not g165(n227, xenc106);
not g166(n222, n332);
not g167(n248, n267);
nand g168(n306, n308, xenc71);
nand g169(n308, add1_i[30], xenc64);
nand g170(n309, add2_i[30], n310);
or g171(n310, xenc64, add1_i[30]);
or g172(n325, add2_i[0], add1_i[0]);
or g173(n342, add2_i[26], add1_i[26]);
nand g174(n286, n288, n289);
nand g175(n289, xenc28, n283);
nand g176(n337, xenc87, xenc82);
nand g177(n345, add2_i[27], add1_i[27]);
nand g178(n346, xenc96, xenc17);
nand g179(n347, n348, xenc46);
nand g180(n348, add2_i[26], add1_i[26]);
nand g181(n294, n296, n297);
nand g182(n296, add2_i[3], add1_i[3]);
nand g183(n297, n298, xenc105);
nand g184(n298, xenc91, n301);
nand g185(n300, add2_i[2], add1_i[2]);
nand g186(n301, n302, xenc98);
not g187(n252, n279);
nand g188(n302, xenc29, n323);
nand g189(n322, add1_i[1], xenc33);
nand g190(n323, add2_i[1], n324);
or g191(n324, xenc33, add1_i[1]);
not g192(n219, add1_i[25]);
not g193(n253, add2_i[25]);
xnor g194(result_o[31], xenc103, xenc92);
xnor g195(n307, add1_i[31], add2_i[31]);
and g196(n315, n335, xenc114);
nand g197(n335, add2_i[28], add1_i[28]);
nand g198(n336, n337, n331);
nand g199(n311, xenc21, n313);
nand g200(n312, add2_i[29], add1_i[29]);
or g201(n313, xenc79, n315);
nand g202(xenc95, n303, n304);
nand g203(n303, add1_i[31], xenc92);
nand g204(n304, add2_i[31], xenc76);
or g205(n305, xenc92, add1_i[31]);
nor g206(n465, add2_i[10], add1_i[10]);
nor g207(n463, add2_i[11], add1_i[11]);
nor g208(n464, add2_i[12], add1_i[12]);
nor g209(n278, add2_i[3], add1_i[3]);
nor g210(n489, add2_i[9], add1_i[9]);
nor g211(n279, add2_i[2], add1_i[2]);
nor g212(n490, add2_i[8], add1_i[8]);
nor g213(n267, n281, n282);
and g214(n282, add1_i[3], xenc60, add2_i[3]);
nor g215(n314, add2_i[29], add1_i[29]);
nand g216(n408, add2_i[14], add1_i[14]);
nand g217(n384, add2_i[17], add1_i[17]);
nand g218(n360, add2_i[20], add1_i[20]);
nand g219(n332, add2_i[23], add1_i[23]);
or g220(n331, add2_i[28], add1_i[28]);
or g221(n440, add2_i[14], add1_i[14]);
or g222(n418, add2_i[17], add1_i[17]);
or g223(n393, add2_i[20], add1_i[20]);
or g224(n369, add2_i[23], add1_i[23]);
or g225(n284, add2_i[6], add1_i[6]);
or g226(n283, add2_i[5], add1_i[5]);
or g227(n266, add2_i[7], add1_i[7]);
nand g228(n484, xenc25, xenc75);
nand g229(n486, n244, n281);
nand g230(n446, xenc5, xenc123);
nand g231(n448, n238, n440);
nand g232(n424, n384, n426);
nand g233(n426, n233, n418);
nand g234(n414, xenc81, n416);
nand g235(n416, n406, xenc10);
nand g236(n399, xenc106, n401);
nand g237(n401, xenc69, xenc120);
nand g238(n389, xenc20, n391);
nand g239(n391, xenc88, xenc52);
nand g240(n375, n332, xenc72);
nand g241(n377, n223, n369);
nand g242(n365, xenc44, xenc1);
nand g243(n367, n358, n225);
nand g244(n351, n348, n353);
nand g245(n353, n218, xenc15);
nand g246(n338, n217, n340);
not g247(n217, n337);
nand g248(n262, xenc49, n265);
nand g249(n265, n266, xenc54, n248);
nand g250(n459, n439, xenc34);
nand g251(n461, n454, xenc14);
nand g252(n273, n247, n275);
nand g253(n275, add2_i[1], add1_i[1], n276, xenc60);
nand g254(n428, n427, n430);
nand g255(n430, xenc65, n431, n241, xenc32);
nand g256(n403, xenc85, n405);
nand g257(n405, xenc107, n406, xenc59, n394);
nand g258(n379, n378, xenc110);
nand g259(n381, n232, xenc88, xenc77, n370);
nand g260(n355, n354, n357);
nand g261(n357, n227, n358, n359, n344);
nand g262(n326, n320, n328);
nand g263(n328, xenc99, xenc101, xenc24, n331);
nand g264(n450, xenc2, xenc112);
nand g265(n452, n453, n454, n245, n441);
xnor g266(n479, add1_i[11], add2_i[11]);
nor g267(n480, xenc50, n476);
nor g268(n481, xenc117, n483, n465);
xnor g269(n471, add1_i[12], add2_i[12]);
nor g270(n472, n473, xenc65);
nor g271(n473, n463, xenc89);
xnor g272(n316, add1_i[30], add2_i[30]);
nor g273(n317, n318, n319);
and g274(n319, add1_i[29], add2_i[29]);
nand g275(n272, n267, n280);
nand g276(n280, add2_i[2], add1_i[2], xenc60, xenc105);
nand g277(n270, add2_i[7], add1_i[7]);
nand g278(n292, add2_i[4], add1_i[4]);
nand g279(n288, add2_i[5], add1_i[5]);
nand g280(n468, add2_i[11], add1_i[11]);
and g281(n458, add1_i[9], add2_i[9]);
and g282(n435, add2_i[12], add1_i[12]);
or g283(n285, add2_i[4], add1_i[4]);
and g284(n453, add2_i[8], add1_i[8]);
or g285(n343, add2_i[27], add1_i[27]);
nand g286(n477, add2_i[6], add1_i[6]);
not g287(n239, add1_i[13]);
not g288(n234, add1_i[16]);
not g289(n236, add1_i[15]);
not g290(n229, add1_i[19]);
not g291(n231, add1_i[18]);
not g292(n224, add1_i[22]);
not g293(n226, add1_i[21]);
not g294(n221, add1_i[24]);
nand g295(n470, add2_i[10], add1_i[10]);
not g296(n261, add2_i[13]);
not g297(n259, add2_i[16]);
not g298(n260, add2_i[15]);
not g299(n257, add2_i[19]);
not g300(n258, add2_i[18]);
not g301(n255, add2_i[22]);
not g302(n256, add2_i[21]);
not g303(n254, add2_i[24]);
nand g304(n436, n417, xenc116);
nand g305(n438, n431, n240);
nand g306(n268, xenc4, xenc22);
nand g307(n271, n272, n266);
nand g308(result_o[0], xenc33, n493);
nand g309(n493, add2_i[0], add1_i[0]);
or g310(xenc0, n457, keyinput0);
or g311(xenc1, n367, keyinput1);
and g312(xenc2, n449, keyinput2);
or g313(xenc3, n411, keyinput3);
and g314(xenc4, n270, keyinput4);
and g315(xenc5, n408, keyinput5);
or g316(xenc6, n470, keyinput6);
or g317(xenc7, n254, keyinput7);
or g318(result_o[24], xenc8, keyinput8);
or g319(result_o[26], xenc9, keyinput9);
or g320(xenc10, n235, keyinput10);
or g321(xenc11, n333, keyinput11);
and g322(xenc12, n269, keyinput12);
and g323(xenc13, n413, keyinput13);
or g324(xenc14, n243, keyinput14);
and g325(xenc15, n342, keyinput15);
or g326(xenc16, n273, keyinput16);
or g327(xenc17, n343, keyinput17);
and g328(xenc18, n420, keyinput18);
or g329(xenc19, n268, keyinput19);
and g330(xenc20, n368, keyinput20);
and g331(xenc21, n312, keyinput21);
or g332(xenc22, n271, keyinput22);
and g333(xenc23, n443, keyinput23);
or g334(xenc24, n330, keyinput24);
and g335(xenc25, n462, keyinput25);
or g336(xenc26, n491, keyinput26);
and g337(result_o[19], xenc27, keyinput27);
and g338(xenc28, n290, keyinput28);
and g339(xenc29, n322, keyinput29);
or g340(xenc30, n385, keyinput30);
or g341(xenc31, n257, keyinput31);
or g342(xenc32, n419, keyinput32);
or g343(xenc33, n325, keyinput33);
or g344(xenc34, n461, keyinput34);
or g345(xenc35, n326, keyinput35);
and g346(xenc36, n455, keyinput36);
and g347(result_o[3], xenc37, keyinput37);
and g348(xenc38, n397, keyinput38);
or g349(xenc39, n471, keyinput39);
or g350(xenc40, n316, keyinput40);
or g351(xenc41, n285, keyinput41);
and g352(xenc42, n460, keyinput42);
and g353(xenc43, n355, keyinput43);
or g354(xenc44, n341, keyinput44);
or g355(xenc45, n490, keyinput45);
and g356(xenc46, n349, keyinput46);
or g357(xenc47, n388, keyinput47);
and g358(xenc48, n224, keyinput48);
and g359(xenc49, n264, keyinput49);
and g360(xenc50, n481, keyinput50);
and g361(xenc51, n459, keyinput51);
or g362(xenc52, n230, keyinput52);
or g363(xenc53, n338, keyinput53);
or g364(xenc54, n246, keyinput54);
and g365(xenc55, n446, keyinput55);
and g366(xenc56, n442, keyinput56);
and g367(xenc57, n414, keyinput57);
and g368(xenc58, n236, keyinput58);
and g369(xenc59, n407, keyinput59);
and g370(xenc60, n277, keyinput60);
and g371(xenc61, n327, keyinput61);
and g372(xenc62, n376, keyinput62);
and g373(xenc63, n364, keyinput63);
or g374(xenc64, n311, keyinput64);
or g375(xenc65, n242, keyinput65);
or g376(xenc66, n286, keyinput66);
or g377(xenc67, n256, keyinput67);
or g378(xenc68, n373, keyinput68);
and g379(xenc69, n228, keyinput69);
and g380(result_o[14], xenc70, keyinput70);
or g381(xenc71, n309, keyinput71);
or g382(xenc72, n377, keyinput72);
and g383(xenc73, n400, keyinput73);
or g384(xenc74, n435, keyinput74);
or g385(xenc75, n486, keyinput75);
or g386(xenc76, n305, keyinput76);
or g387(xenc77, n383, keyinput77);
and g388(xenc78, n260, keyinput78);
and g389(xenc79, n314, keyinput79);
and g390(xenc80, n292, keyinput80);
and g391(xenc81, n392, keyinput81);
and g392(xenc82, n346, keyinput82);
or g393(xenc83, n239, keyinput83);
and g394(result_o[13], xenc84, keyinput84);
or g395(xenc85, n402, keyinput85);
or g396(result_o[27], xenc86, keyinput86);
and g397(xenc87, n345, keyinput87);
or g398(xenc88, n382, keyinput88);
or g399(xenc89, n474, keyinput89);
and g400(result_o[1], xenc90, keyinput90);
and g401(xenc91, n300, keyinput91);
or g402(xenc92, n306, keyinput92);
and g403(result_o[15], xenc93, keyinput93);
and g404(xenc94, n444, keyinput94);
or g405(result_o[32], xenc95, keyinput95);
or g406(xenc96, n347, keyinput96);
or g407(xenc97, n399, keyinput97);
and g408(xenc98, n252, keyinput98);
or g409(xenc99, n222, keyinput99);
or g410(result_o[8], xenc100, keyinput100);
or g411(xenc101, n329, keyinput101);
and g412(xenc102, n299, keyinput102);
or g413(xenc103, n307, keyinput103);
or g414(xenc104, n429, keyinput104);
or g415(xenc105, n251, keyinput105);
and g416(xenc106, n360, keyinput106);
or g417(xenc107, n237, keyinput107);
and g418(result_o[12], xenc108, keyinput108);
and g419(xenc109, n484, keyinput109);
or g420(xenc110, n381, keyinput110);
and g421(xenc111, n258, keyinput111);
and g422(xenc112, n452, keyinput112);
or g423(xenc113, n356, keyinput113);
or g424(xenc114, n336, keyinput114);
and g425(xenc115, n432, keyinput115);
or g426(xenc116, n438, keyinput116);
and g427(xenc117, n478, keyinput117);
and g428(xenc118, n428, keyinput118);
and g429(result_o[5], xenc119, keyinput119);
and g430(xenc120, n393, keyinput120);
or g431(xenc121, n451, keyinput121);
and g432(xenc122, n403, keyinput122);
or g433(xenc123, n448, keyinput123);
or g434(xenc124, n467, keyinput124);
and g435(xenc125, n250, keyinput125);
and g436(xenc126, n409, keyinput126);
or g437(result_o[23], xenc127, keyinput127);
endmodule
