library verilog;
use verilog.vl_types.all;
entity ripple_carry_adder32_tb is
end ripple_carry_adder32_tb;
