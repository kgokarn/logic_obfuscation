// Verilog File 
module carry_lookahead_adder32_xor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n659, xenc93, xenc52, n660, xenc99, xenc0, xenc41, n664, xenc111, 
n666, xenc8, n668, n669, xenc96, xenc88, xenc51, n679, n684, n685, 
xenc28, n690, n691, xenc35, xenc1, xenc27, xenc25, n701, n872, xenc45, 
xenc106, n711, xenc92, n721, xenc44, xenc127, xenc43, xenc119, n731, n736, 
n737, xenc67, xenc22, xenc29, xenc75, n743, n752, xenc49, n753, xenc71, 
n763, xenc82, n772, xenc4, xenc31, n773, xenc48, xenc117, n783, n830, 
n826, n832, n828, n836, n838, n834, n814, n815, n665, xenc59, 
n802, n816, n827, xenc24, n817, xenc17, n889, xenc33, n769, n818, 
n819, n833, xenc91, n820, n821, n839, n822, n749, n831, n823, 
xenc114, n829, xenc80, xenc55, n824, n825, n770, xenc15, n785, n864, 
n788, n750, xenc95, n740, n835, n888, n890, n875, xenc61, n837, 
n775, xenc13, xenc109, n745, xenc123, xenc97, n840, n841, xenc87, xenc9, 
n842, n683, n843, n715, n844, xenc65, n655, xenc98, xenc58, n845, 
n846, n847, n729, n799, xenc11, n849, n876, n871, n848, xenc50, 
xenc126, xenc72, xenc32, n891, xenc16, n850, n860, xenc38, n851, n852, 
xenc63, xenc37, n853, xenc39, xenc103, n854, n757, xenc56, n726, n855, 
xenc120, xenc46, n856, xenc124, xenc20, xenc115, n857, xenc78, xenc7, n858, 
n656, xenc18, xenc113, xenc3, n859, n861, n717, xenc76, n714, xenc104, 
xenc68, n862, n863, n865, n780, xenc53, n866, xenc116, n707, xenc47, 
xenc81, n867, n868, n869, n870, n708, n873, xenc57, n874, xenc30, 
xenc112, n703, n880, n877, xenc110, n722, n879, xenc101, n878, n881, 
xenc89, n724, n882, xenc85, n725, n806, n805, xenc86, xenc14, n792, 
xenc2, xenc36, n883, n884, n662, xenc70, n885, xenc26, xenc23, n795, 
n887, xenc5, n886, n813, n798, n663, xenc42, n676, xenc69, n688, 
n687, xenc34, n747, xenc74, n767, xenc83, xenc54, n765, xenc100, n755, 
n812, n811, n810, n658, xenc118, n705, n670, n671, xenc64, n698, 
n695, n719, n718, n727, n760, n787, xenc66, n794, n804, n807, 
n809, n728, xenc21, xenc19, n702, n700, xenc125, n754, xenc121, n808, 
n732, xenc90, n730, n734, n733, n774, xenc108, n791, xenc12, n675, 
n677, n689, n739, n759, n761, n779, xenc77, xenc40, n673, xenc73, 
n735, xenc107, n777, n680, n681, n678, n682, xenc10, n693, n694, 
xenc94, n723, n720, xenc84, n742, xenc102, xenc6, n762, n784, n782, 
xenc60, n803, xenc105, xenc62, xenc122, n672, n692, n697, n699, n712, 
n744, n764, n790, n793, xenc79;

xor g0(xenc52, n659, xenc93);
xor g1(n660, add2_i[8], add1_i[8]);
xor g2(xenc41, xenc99, xenc0);
xor g3(n664, add2_i[6], add1_i[6]);
xor g4(xenc8, xenc111, n666);
xor g5(n666, add2_i[5], add1_i[5]);
xor g6(result_o[3], n668, n669);
xor g7(n669, add2_i[3], add1_i[3]);
xor g8(xenc51, xenc96, xenc88);
xor g9(n679, add2_i[30], add1_i[30]);
xor g10(xenc28, n684, n685);
xor g11(n685, add2_i[2], add1_i[2]);
xor g12(xenc35, n690, n691);
xor g13(n691, add2_i[28], add1_i[28]);
xor g14(xenc25, xenc1, xenc27);
xor g15(n701, add2_i[26], add1_i[26]);
xor g16(xenc106, n872, xenc45);
xor g17(n711, add2_i[24], add1_i[24]);
xor g18(xenc44, xenc92, n721);
xor g19(n721, add2_i[22], add1_i[22]);
xor g20(xenc119, xenc127, xenc43);
xor g21(n731, add2_i[20], add1_i[20]);
xor g22(xenc67, n736, n737);
xor g23(n737, add2_i[1], add1_i[1]);
xor g24(xenc75, xenc22, xenc29);
xor g25(n743, add2_i[18], add1_i[18]);
xor g26(result_o[16], n752, xenc49);
xor g27(n753, add2_i[16], add1_i[16]);
xor g28(xenc82, xenc71, n763);
xor g29(n763, add2_i[14], add1_i[14]);
xor g30(xenc31, n772, xenc4);
xor g31(n773, add2_i[12], add1_i[12]);
xor g32(result_o[10], xenc48, xenc117);
xor g33(n783, add2_i[10], add1_i[10]);
or g34(n736, add2_i[0], add1_i[0]);
not g35(n830, add2_i[8]);
not g36(n826, add2_i[12]);
not g37(n832, add2_i[16]);
not g38(n828, add2_i[9]);
not g39(n836, add2_i[11]);
not g40(n838, add2_i[17]);
not g41(n834, add2_i[18]);
nand g42(n665, n814, n815);
nand g43(n814, add1_i[4], xenc59);
nand g44(n815, add2_i[4], n802);
or g45(n816, add2_i[0], add1_i[1]);
or g46(n817, n827, xenc24);
and g47(n889, n817, xenc17);
and g48(n818, xenc33, n769);
not g49(n819, add1_i[13]);
or g50(n820, n833, xenc91);
and g51(n839, n820, n821);
and g52(n821, n822, n749);
not g53(n822, add1_i[17]);
or g54(n823, n831, n830);
and g55(n829, n823, xenc114);
and g56(n824, xenc80, xenc55);
not g57(n825, add1_i[9]);
or g58(n770, xenc24, n827);
nor g59(n827, n772, add1_i[12]);
or g60(n785, n829, xenc15);
not g61(n864, add2_i[10]);
or g62(n788, n830, n831);
nor g63(n831, n659, add1_i[8]);
or g64(n750, xenc91, n833);
nor g65(n833, n752, add1_i[16]);
or g66(n740, n834, xenc95);
nor g67(n835, xenc22, add1_i[18]);
not g68(n888, add2_i[13]);
not g69(n890, add2_i[15]);
not g70(n875, add2_i[25]);
or g71(n775, xenc61, n837);
nor g72(n837, xenc13, add1_i[11]);
or g73(n745, xenc109, n839);
xor g74(result_o[31], xenc123, xenc97);
xor g75(n840, add1_i[31], add2_i[31]);
xor g76(xenc9, n841, xenc87);
xor g77(n841, add1_i[27], add2_i[27]);
xor g78(result_o[29], n842, n683);
xor g79(n842, add1_i[29], add2_i[29]);
xor g80(result_o[23], n843, n715);
xor g81(n843, add1_i[23], add2_i[23]);
xor g82(result_o[25], n844, xenc65);
xor g83(n844, add1_i[25], add2_i[25]);
not g84(n655, add1_i[4]);
nor g85(n845, xenc98, xenc58);
and g86(n846, add1_i[5], n802, add2_i[4]);
and g87(n847, add1_i[5], xenc59, add1_i[4]);
or g88(n729, xenc127, add1_i[20]);
or g89(n799, xenc111, add1_i[5]);
nor g90(n876, xenc11, n849);
and g91(n848, n871, add2_i[24]);
nand g92(n849, xenc50, xenc126);
nor g93(n891, xenc72, xenc32);
and g94(n850, xenc16, add2_i[14]);
nand g95(n851, n860, xenc38);
xor g96(xenc37, n852, xenc63);
xor g97(n852, add1_i[17], add2_i[17]);
xor g98(xenc103, n853, xenc39);
xor g99(n853, add1_i[19], add2_i[19]);
xor g100(xenc56, n854, n757);
xor g101(n854, add1_i[15], add2_i[15]);
xnor g102(n726, add1_i[21], add2_i[21]);
xor g103(xenc46, n855, xenc120);
xor g104(n855, add1_i[13], add2_i[13]);
xor g105(result_o[9], n856, xenc124);
xor g106(n856, add1_i[9], add2_i[9]);
xor g107(xenc115, xenc20, xenc13);
xor g108(n857, add1_i[11], add2_i[11]);
xor g109(result_o[7], xenc78, xenc7);
xor g110(n858, add1_i[7], add2_i[7]);
xor g111(xenc113, n656, xenc18);
xor g112(n859, add2_i[4], xenc3);
not g113(n860, add1_i[15]);
not g114(n861, add1_i[25]);
nand g115(n714, n717, xenc76);
and g116(n862, xenc104, xenc68);
not g117(n863, add1_i[23]);
or g118(n780, n865, n864);
nor g119(n865, xenc48, add1_i[10]);
nand g120(n866, n714, xenc53);
and g121(n707, n866, xenc116);
or g122(n867, xenc47, xenc81);
not g123(n868, add1_i[24]);
and g124(n869, add2_i[23], add1_i[24]);
nand g125(n870, add2_i[23], n714);
nand g126(n708, n871, add2_i[24]);
nand g127(n871, n873, xenc57);
nand g128(n872, xenc81, n870);
nand g129(n873, n714, add2_i[23]);
and g130(n874, xenc47, xenc81);
or g131(n703, xenc30, xenc112);
nand g132(n877, n729, n880);
and g133(n722, n877, xenc110);
or g134(n878, n879, xenc101);
not g135(n879, add1_i[21]);
and g136(n880, add2_i[20], add1_i[21]);
nand g137(n881, n729, add2_i[20]);
nand g138(n724, n881, xenc89);
and g139(n882, n879, xenc101);
nand g140(n725, xenc101, xenc85);
nand g141(n805, add2_i[3], n806);
nand g142(n792, xenc86, xenc14);
and g143(n883, xenc2, xenc36);
not g144(n884, add1_i[7]);
nand g145(n662, xenc14, xenc2);
nand g146(n885, xenc70, add2_i[5]);
nand g147(n795, xenc26, xenc23);
and g148(n886, n887, xenc5);
not g149(n887, add1_i[6]);
nand g150(n813, add2_i[0], add1_i[0]);
nand g151(n663, n798, xenc5);
nand g152(n676, add2_i[30], xenc42);
nand g153(n798, xenc70, add2_i[5]);
nand g154(n688, add2_i[28], xenc69);
nand g155(n683, n687, n688);
nand g156(n747, n749, xenc34);
nand g157(n767, n769, xenc74);
or g158(n765, xenc83, xenc54);
or g159(n755, xenc100, n891);
nand g160(n811, add2_i[1], n812);
nand g161(n684, n810, n811);
nand g162(n658, xenc55, n788);
nand g163(n705, xenc126, xenc118);
nand g164(result_o[32], n670, n671);
nand g165(n695, xenc64, n698);
nand g166(n718, add2_i[22], n719);
nand g167(n727, add1_i[20], xenc127);
nand g168(n760, add2_i[14], xenc16);
nand g169(n769, add1_i[12], n772);
nand g170(n787, add1_i[8], n659);
nand g171(n794, add2_i[6], xenc66);
nand g172(n804, add1_i[3], n668);
or g173(n806, n668, add1_i[3]);
nand g174(n807, add1_i[2], n684);
or g175(n809, n684, add1_i[2]);
nand g176(n728, add2_i[20], n729);
nand g177(n671, add2_i[31], xenc21);
nand g178(n698, add2_i[26], xenc19);
nand g179(n700, n703, n702);
nand g180(n752, xenc125, n754);
nand g181(n668, xenc121, n808);
nand g182(n808, add2_i[2], n809);
nand g183(n730, n732, xenc90);
nand g184(n733, add2_i[19], n734);
nand g185(n772, n774, n775);
nand g186(n659, xenc108, n791);
nand g187(n791, xenc12, add2_i[7]);
nand g188(n675, add1_i[30], xenc96);
or g189(n677, xenc96, add1_i[30]);
nand g190(n687, add1_i[28], n690);
or g191(n689, n690, add1_i[28]);
nand g192(n717, add1_i[22], xenc92);
or g193(n719, xenc92, add1_i[22]);
nand g194(n739, add1_i[18], xenc22);
nand g195(n759, add1_i[14], xenc71);
or g196(n761, xenc71, add1_i[14]);
nand g197(n779, add1_i[10], xenc48);
nand g198(n673, xenc77, xenc40);
nand g199(n715, n717, xenc104);
nand g200(n735, xenc73, n740);
nand g201(n757, xenc38, xenc107);
nand g202(n777, n780, n779);
nand g203(n802, n656, xenc3);
nand g204(n678, n680, n681);
nand g205(n681, add2_i[29], n682);
nand g206(n690, xenc10, n693);
nand g207(n693, add2_i[27], n694);
nand g208(n720, xenc94, n723);
nand g209(n723, n724, add2_i[21]);
nand g210(n742, xenc84, n745);
nand g211(n762, xenc102, xenc6);
nand g212(n782, n784, n785);
nand g213(n803, n805, xenc60);
nand g214(xenc105, n736, n813);
xnor g215(result_o[21], xenc62, xenc122);
nand g216(n670, add1_i[31], xenc97);
or g217(n672, xenc97, add1_i[31]);
nand g218(n680, add1_i[29], n683);
or g219(n682, n683, add1_i[29]);
nand g220(n692, add1_i[27], xenc87);
or g221(n694, xenc87, add1_i[27]);
nand g222(n697, add1_i[26], xenc1);
or g223(n699, xenc1, add1_i[26]);
nand g224(n702, add1_i[25], xenc65);
nand g225(n712, add1_i[23], n715);
nand g226(n732, add1_i[19], xenc39);
or g227(n734, xenc39, add1_i[19]);
nand g228(n744, add1_i[17], xenc63);
nand g229(n749, add1_i[16], n752);
nand g230(n754, add1_i[15], n757);
nand g231(n764, add1_i[13], xenc120);
nand g232(n774, add1_i[11], xenc13);
nand g233(n784, add1_i[9], xenc124);
nand g234(n790, add1_i[7], xenc7);
nand g235(n793, add1_i[6], xenc99);
not g236(n656, xenc59);
nand g237(n810, add1_i[1], n736);
or g238(n812, xenc79, add1_i[0]);
xor g239(xenc0, n664, keyinput0);
xnor g240(xenc1, n700, keyinput1);
xnor g241(xenc2, n794, keyinput2);
xnor g242(xenc3, n655, keyinput3);
xnor g243(xenc4, n773, keyinput4);
xor g244(xenc5, n845, keyinput5);
xor g245(xenc6, n765, keyinput6);
xor g246(xenc7, n662, keyinput7);
xor g247(result_o[5], xenc8, keyinput8);
xnor g248(result_o[27], xenc9, keyinput9);
xor g249(xenc10, n692, keyinput10);
xor g250(xenc11, n848, keyinput11);
xor g251(xenc12, n792, keyinput12);
xor g252(xenc13, n777, keyinput13);
xor g253(xenc14, n793, keyinput14);
xor g254(xenc15, n828, keyinput15);
xor g255(xenc16, n761, keyinput16);
xor g256(xenc17, n818, keyinput17);
xnor g257(xenc18, n859, keyinput18);
xnor g258(xenc19, n699, keyinput19);
xor g259(xenc20, n857, keyinput20);
xor g260(xenc21, n672, keyinput21);
xnor g261(xenc22, n742, keyinput22);
xnor g262(xenc23, n886, keyinput23);
xor g263(xenc24, n826, keyinput24);
xnor g264(result_o[26], xenc25, keyinput25);
xnor g265(xenc26, n885, keyinput26);
xor g266(xenc27, n701, keyinput27);
xnor g267(result_o[2], xenc28, keyinput28);
xor g268(xenc29, n743, keyinput29);
xnor g269(xenc30, n876, keyinput30);
xor g270(result_o[12], xenc31, keyinput31);
xnor g271(xenc32, n851, keyinput32);
xnor g272(xenc33, n819, keyinput33);
xor g273(xenc34, n750, keyinput34);
xnor g274(result_o[28], xenc35, keyinput35);
xnor g275(xenc36, n884, keyinput36);
xor g276(result_o[17], xenc37, keyinput37);
xor g277(xenc38, n759, keyinput38);
xor g278(xenc39, n735, keyinput39);
xor g279(xenc40, n676, keyinput40);
xnor g280(result_o[6], xenc41, keyinput41);
xnor g281(xenc42, n677, keyinput42);
xor g282(xenc43, n731, keyinput43);
xor g283(result_o[22], xenc44, keyinput44);
xor g284(xenc45, n711, keyinput45);
xnor g285(result_o[13], xenc46, keyinput46);
xnor g286(xenc47, n868, keyinput47);
xnor g287(xenc48, n782, keyinput48);
xnor g288(xenc49, n753, keyinput49);
xor g289(xenc50, n861, keyinput50);
xor g290(result_o[30], xenc51, keyinput51);
xor g291(result_o[8], xenc52, keyinput52);
xor g292(xenc53, n869, keyinput53);
xnor g293(xenc54, n889, keyinput54);
xnor g294(xenc55, n787, keyinput55);
xnor g295(result_o[15], xenc56, keyinput56);
xnor g296(xenc57, n874, keyinput57);
xnor g297(xenc58, n847, keyinput58);
xnor g298(xenc59, n803, keyinput59);
xor g299(xenc60, n804, keyinput60);
xnor g300(xenc61, n836, keyinput61);
xor g301(xenc62, n726, keyinput62);
xor g302(xenc63, n747, keyinput63);
xnor g303(xenc64, n697, keyinput64);
xnor g304(xenc65, n705, keyinput65);
xnor g305(xenc66, n795, keyinput66);
xnor g306(result_o[1], xenc67, keyinput67);
xor g307(xenc68, n863, keyinput68);
xor g308(xenc69, n689, keyinput69);
xor g309(xenc70, n799, keyinput70);
xor g310(xenc71, n762, keyinput71);
xnor g311(xenc72, n850, keyinput72);
xnor g312(xenc73, n739, keyinput73);
xnor g313(xenc74, n770, keyinput74);
xor g314(result_o[18], xenc75, keyinput75);
xor g315(xenc76, n862, keyinput76);
xnor g316(xenc77, n675, keyinput77);
xnor g317(xenc78, n858, keyinput78);
xnor g318(xenc79, n816, keyinput79);
xnor g319(xenc80, n825, keyinput80);
xor g320(xenc81, n712, keyinput81);
xor g321(result_o[14], xenc82, keyinput82);
xor g322(xenc83, n888, keyinput83);
xnor g323(xenc84, n744, keyinput84);
xor g324(xenc85, n728, keyinput85);
xnor g325(xenc86, n883, keyinput86);
xnor g326(xenc87, n695, keyinput87);
xor g327(xenc88, n679, keyinput88);
xnor g328(xenc89, n882, keyinput89);
xnor g329(xenc90, n733, keyinput90);
xor g330(xenc91, n832, keyinput91);
xnor g331(xenc92, n720, keyinput92);
xor g332(xenc93, n660, keyinput93);
xnor g333(xenc94, n722, keyinput94);
xnor g334(xenc95, n835, keyinput95);
xnor g335(xenc96, n678, keyinput96);
xnor g336(xenc97, n673, keyinput97);
xor g337(xenc98, n846, keyinput98);
xor g338(xenc99, n663, keyinput99);
xnor g339(xenc100, n890, keyinput100);
xnor g340(xenc101, n727, keyinput101);
xnor g341(xenc102, n764, keyinput102);
xnor g342(result_o[19], xenc103, keyinput103);
xnor g343(xenc104, n718, keyinput104);
xnor g344(result_o[0], xenc105, keyinput105);
xor g345(result_o[24], xenc106, keyinput106);
xnor g346(xenc107, n760, keyinput107);
xnor g347(xenc108, n790, keyinput108);
xor g348(xenc109, n838, keyinput109);
xnor g349(xenc110, n878, keyinput110);
xnor g350(xenc111, n665, keyinput111);
xnor g351(xenc112, n875, keyinput112);
xor g352(result_o[4], xenc113, keyinput113);
xnor g353(xenc114, n824, keyinput114);
xor g354(result_o[11], xenc115, keyinput115);
xor g355(xenc116, n867, keyinput116);
xnor g356(xenc117, n783, keyinput117);
xor g357(xenc118, n708, keyinput118);
xnor g358(result_o[20], xenc119, keyinput119);
xnor g359(xenc120, n767, keyinput120);
xnor g360(xenc121, n807, keyinput121);
xor g361(xenc122, n725, keyinput122);
xnor g362(xenc123, n840, keyinput123);
xor g363(xenc124, n658, keyinput124);
xnor g364(xenc125, n755, keyinput125);
xnor g365(xenc126, n707, keyinput126);
xor g366(xenc127, n730, keyinput127);
endmodule
