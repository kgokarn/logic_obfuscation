module xnor_based_carry_lookahead_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141;

  xor U132 ( result_o[9], n64, n65);
  xor U133 ( n65, add2_i[9], add1_i[9]);
  xor U134 ( result_o[8], n66, n67);
  xor U135 ( n67, add2_i[8], add1_i[8]);
  xor U136 ( result_o[7], n68, n69);
  xor U137 ( n69, add2_i[7], add1_i[7]);
  xor U138 ( result_o[6], n70, n71);
  xor U139 ( n71, add2_i[6], add1_i[6]);
  xor U140 ( result_o[5], n72, n73);
  xor U141 ( n73, add2_i[5], add1_i[5]);
  xor U142 ( result_o[4], n74, n75);
  xor U143 ( n75, add2_i[4], add1_i[4]);
  xor U146 ( n81, add2_i[1], add1_i[1]);
  xor U147 ( result_o[15], n85, n86);
  xor U148 ( n86, add2_i[15], add1_i[15]);
  xor U149 ( result_o[14], n90, n91);
  xor U150 ( n91, add2_i[14], add1_i[14]);
  xor U151 ( result_o[13], n95, n96);
  xor U152 ( n96, add2_i[13], add1_i[13]);
  xor U153 ( result_o[12], n100, n101);
  xor U154 ( n101, add2_i[12], add1_i[12]);
  xor U155 ( result_o[11], n105, n106);
  xor U156 ( n106, add2_i[11], add1_i[11]);
  xor U157 ( result_o[10], n110, n111);
  xor U158 ( n111, add2_i[10], add1_i[10]);
  not U159 ( n63, n80);
  nor U160 ( n80, add2_i[0], add1_i[0]);
  nand U161 ( n72, n127, n128);
  nand U162 ( n127, add1_i[4], n74);
  nand U163 ( n128, add2_i[4], n129);
  or U164 ( n129, n74, add1_i[4]);
  nand U165 ( n95, n97, n98);
  nand U166 ( n97, add1_i[12], n100);
  nand U167 ( n98, add2_i[12], n99);
  or U168 ( n99, n100, add1_i[12]);
  nand U169 ( n90, n92, n93);
  nand U170 ( n92, add1_i[13], n95);
  nand U171 ( n93, add2_i[13], n94);
  or U172 ( n94, n95, add1_i[13]);
  nand U173 ( n85, n87, n88);
  nand U174 ( n87, add1_i[14], n90);
  nand U175 ( n88, add2_i[14], n89);
  or U176 ( n89, n90, add1_i[14]);
  nand U177 ( n79, n136, n137);
  nand U178 ( n136, add1_i[1], n63);
  nand U179 ( n137, add2_i[1], n138);
  or U180 ( n138, n63, add1_i[1]);
  nand U181 ( n77, n133, n134);
  nand U182 ( n133, add1_i[2], n79);
  nand U183 ( n134, add2_i[2], n135);
  or U184 ( n135, n79, add1_i[2]);
  nand U185 ( n74, n130, n131);
  nand U186 ( n130, add1_i[3], n77);
  nand U187 ( n131, add2_i[3], n132);
  or U188 ( n132, n77, add1_i[3]);
  nand U189 ( n70, n124, n125);
  nand U190 ( n124, add1_i[5], n72);
  nand U191 ( n125, add2_i[5], n126);
  or U192 ( n126, n72, add1_i[5]);
  nand U193 ( n68, n121, n122);
  nand U194 ( n121, add1_i[6], n70);
  nand U195 ( n122, add2_i[6], n123);
  or U196 ( n123, n70, add1_i[6]);
  nand U197 ( n66, n118, n119);
  nand U198 ( n118, add1_i[7], n68);
  nand U199 ( n119, add2_i[7], n120);
  or U200 ( n120, n68, add1_i[7]);
  nand U201 ( n64, n115, n116);
  nand U202 ( n115, add1_i[8], n66);
  nand U203 ( n116, add2_i[8], n117);
  or U204 ( n117, n66, add1_i[8]);
  nand U205 ( n110, n112, n113);
  nand U206 ( n112, add1_i[9], n64);
  nand U207 ( n113, add2_i[9], n114);
  or U208 ( n114, n64, add1_i[9]);
  nand U209 ( n105, n107, n108);
  nand U210 ( n107, add1_i[10], n110);
  nand U211 ( n108, add2_i[10], n109);
  or U212 ( n109, n110, add1_i[10]);
  nand U213 ( n100, n102, n103);
  nand U214 (n102, add1_i[11], n105);
  nand U215 ( n103, add2_i[11], n104);
  or U216 ( n104, n105, add1_i[11]);
  nand U217 ( result_o[16], n82, n83);
  nand U218 ( n82, add1_i[15], n85);
  nand U219 ( n83, add2_i[15], n84);
  or U220 ( n84, n85, add1_i[15]);
  nor U221 ( result_o[1], n80, n81);
  and U222 ( result_o[2], n79, n140);
  xnor U223 ( n140, add2_i[2], add1_i[2]);
  and U224 ( result_o[3], n77, n141);
  xnor U225 ( n141, add2_i[3], add1_i[3]);
  nand U226 ( result_o[0], n63, n139);
  nand U227 ( n139, add2_i[0], add1_i[0]);
endmodule
