module equal_segmentation_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181;

  xor U84 ( result_o[9], add2_i[9], n76);
  xor U85 ( result_o[8], add2_i[8], add1_i[8]);
  xor U86 ( result_o[7], n77, n78);
  xor U87 ( n78, add2_i[7], add1_i[7]);
  xor U88 ( result_o[6], add2_i[6], n81);
  xor U89 ( n81, n82, add1_i[6]);
  xor U90 ( result_o[5], add2_i[5], n85);
  xor U91 ( n85, n86, add1_i[5]);
  xor U92 ( result_o[4], add2_i[4], n89);
  xor U93 ( n89, n90, add1_i[4]);
  xor U94 ( result_o[3], add2_i[3], n93);
  xor U95 ( n93, n94, add1_i[3]);
  xor U96 ( result_o[31], add2_i[31], n101);
  xor U97 ( n101, n102, add1_i[31]);
  xor U98 ( result_o[30], add2_i[30], n105);
  xor U99 ( n105, n106, add1_i[30]);
  xor U100 ( result_o[2], add2_i[2], n97);
  xor U101 ( n97, n98, add1_i[2]);
  xor U102 ( result_o[29], add2_i[29], n109);
  xor U103 ( n109, n110, add1_i[29]);
  xor U104 ( result_o[28], add2_i[28], n116);
  xor U105 ( n116, n117, add1_i[28]);
  xor U106 ( result_o[27], add2_i[27], n120);
  xor U107 ( n120, n121, add1_i[27]);
  xor U108 ( result_o[26], add2_i[26], n124);
  xor U109 ( n124, n125, add1_i[26]);
  xor U110 ( result_o[25], add2_i[25], n128);
  xor U111 ( result_o[24], add2_i[24], add1_i[24]);
  xor U112 ( result_o[23], n130, n131);
  xor U113 ( n131, add2_i[23], add1_i[23]);
  xor U114 ( result_o[22], add2_i[22], n134);
  xor U115 ( n134, n135, add1_i[22]);
  xor U116 ( result_o[21], add2_i[21], n138);
  xor U117 ( n138, n139, add1_i[21]);
  xor U118 ( result_o[20], add2_i[20], n142);
  xor U119 ( n142, n143, add1_i[20]);
  xor U120 ( result_o[1], add2_i[1], n113);
  xor U121 ( result_o[19], add2_i[19], n146);
  xor U122 ( n146, n147, add1_i[19]);
  xor U123 ( result_o[18], add2_i[18], n151);
  xor U124 ( n151, n152, add1_i[18]);
  xor U125 ( result_o[17], add2_i[17], n155);
  xor U126 ( result_o[16], add2_i[16], add1_i[16]);
  xor U127 ( result_o[15], n157, n158);
  xor U128 ( n158, add2_i[15], add1_i[15]);
  xor U129 ( result_o[14], add2_i[14], n161);
  xor U130 ( n161, n162, add1_i[14]);
  xor U131 ( result_o[13], add2_i[13], n165);
  xor U132 ( n165, n166, add1_i[13]);
  xor U133 ( result_o[12], add2_i[12], n169);
  xor U134 ( n169, n170, add1_i[12]);
  xor U135 ( result_o[11], add2_i[11], n173);
  xor U136 ( n173, n174, add1_i[11]);
  xor U137 ( result_o[10], add2_i[10], n177);
  xor U138 ( n177, n178, add1_i[10]);
  xor U139 ( result_o[0], add2_i[0], add1_i[0]);
  xnor U140 ( n128, n129, add1_i[25]);
  nand U141 ( n129, add2_i[24], add1_i[24]);
  xnor U142 ( n113, n148, add1_i[1]);
  nand U143 ( n148, add2_i[0], add1_i[0]);
  xnor U144 ( n76, n181, add1_i[9]);
  nand U145 ( n181, add2_i[8], add1_i[8]);
  xnor U146 ( n155, n156, add1_i[17]);
  nand U147 ( n156, add2_i[16], add1_i[16]);
  nand U148 ( n77, n79, n80);
  nand U149 ( n79, add1_i[6], n82);
  nand U150 ( n157, n159, n160);
  nand U151 ( n159, add1_i[14], n162);
  nand U152 ( n130, n132, n133);
  nand U153 ( n132, add1_i[22], n135);
  nand U154 ( n121, n122, n123);
  nand U155 ( n122, add1_i[26], n125);
  nand U156 ( n123, add2_i[26], n124);
  nand U157 ( n94, n95, n96);
  nand U158 ( n95, add1_i[2], n98);
  nand U159 ( n96, add2_i[2], n97);
  nand U160 ( n174, n175, n176);
  nand U161 ( n175, add1_i[10], n178);
  nand U162 ( n176, add2_i[10], n177);
  nand U163 ( n147, n149, n150);
  nand U164 ( n149, add1_i[18], n152);
  nand U165 ( n150, add2_i[18], n151);
  nand U166 ( n117, n118, n119);
  nand U167 ( n118, add1_i[27], n121);
  nand U168 ( n119, add2_i[27], n120);
  nand U169 ( n90, n91, n92);
  nand U170 ( n91, add1_i[3], n94);
  nand U171 ( n92, add2_i[3], n93);
  nand U172 ( n170, n171, n172);
  nand U173 ( n171, add1_i[11], n174);
  nand U174 ( n172, add2_i[11], n173);
  nand U175 ( n143, n144, n145);
  nand U176 ( n144, add1_i[19], n147);
  nand U177 ( n145, add2_i[19], n146);
  nand U178 ( n102, n103, n104);
  nand U179 ( n103, add1_i[30], n106);
  nand U180 ( n104, add2_i[30], n105);
  nand U181 ( n110, n114, n115);
  nand U182 ( n114, add1_i[28], n117);
  nand U183 ( n115, add2_i[28], n116);
  nand U184 ( n86, n87, n88);
  nand U185 ( n87, add1_i[4], n90);
  nand U186 ( n88, add2_i[4], n89);
  nand U187 ( n166, n167, n168);
  nand U188 ( n167, add1_i[12], n170);
  nand U189 ( n168, add2_i[12], n169);
  nand U190 ( n139, n140, n141);
  nand U191 ( n140, add1_i[20], n143);
  nand U192 ( n141, add2_i[20], n142);
  nand U193 ( n106, n107, n108);
  nand U194 ( n107, add1_i[29], n110);
  nand U195 ( n108, add2_i[29], n109);
  nand U196 ( n82, n83, n84);
  nand U197 ( n83, add1_i[5], n86);
  nand U198 ( n84, add2_i[5], n85);
  nand U199 ( n162, n163, n164);
  nand U200 ( n163, add1_i[13], n166);
  nand U201 ( n164, add2_i[13], n165);
  nand U202 ( n135, n136, n137);
  nand U203 ( n136, add1_i[21], n139);
  nand U204 ( n137, add2_i[21], n138);
  nand U205 ( n80, add2_i[6], n81);
  nand U206 ( n160, add2_i[14], n161);
  nand U207 ( n133, add2_i[22], n134);
  nand U208 ( n125, n126, n127);
  nand U209 ( n127, add1_i[25], add1_i[24], add2_i[24]);
  nand U210 ( n126, add2_i[25], n128);
  nand U211 ( n98, n111, n112);
  nand U212 ( n112, add1_i[1], add1_i[0], add2_i[0]);
  nand U213 ( n111, add2_i[1], n113);
  nand U214 ( n178, n179, n180);
  nand U215 ( n180, add2_i[8], add1_i[8], add1_i[9]);
  nand U216 ( n179, add2_i[9], n76);
  nand U217 ( n152, n153, n154);
  nand U218 ( n154, add1_i[17], add1_i[16], add2_i[16]);
  nand U219 ( n153, add2_i[17], n155);
  nand U220 ( result_o[32], n99, n100);
  nand U221 ( n99, add1_i[31], n102);
  nand U222 ( n100, add2_i[31], n101);
endmodule
