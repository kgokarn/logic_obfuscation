module broke_array_multiplier8 ( op1_i, op2_i, product_o );
  input [7:0] op1_i, op2_i;
  output [15:0] product_o;
  wire   n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487;

  xor U280 ( product_o[9], n203, n204);
  xor U281 ( n203, n205, n206);
  xor U283 ( product_o[14], n222, n223);
  xor U284 ( product_o[13], n238, n237);
  xor U285 ( n237, n230, n239);
  xor U286 ( n239, n229, n231);
  xor U287 ( n238, n236, n234);
  xor U288 ( product_o[12], n258, n257);
  xor U289 ( n258, n256, n254);
  xor U290 ( product_o[11], n282, n283);
  xor U291 ( n283, n281, n279);
  xor U292 ( n275, n269, n298);
  xor U293 ( n208, n325, n326);
  xor U294 ( n325, n327, n328);
  xor U295 ( n330, n347, n348);
  xor U296 ( n347, n349, n350);
  xor U297 ( n319, n355, n356);
  xor U298 ( n296, n359, n312);
  xor U299 ( n307, n301, n361);
  xor U300 ( n359, n313, n310);
  xor U301 ( n348, n383, n384);
  xor U302 ( n383, n385, n386);
  xor U303 ( n352, n390, n391);
  xor U304 ( n390, n392, n393);
  xor U305 ( n341, n398, n399);
  xor U306 ( n355, n402, n373);
  xor U307 ( n402, n372, n370);
  xor U308 ( n384, n441, n442);
  xor U309 ( n442, n443, n444);
  xor U310 ( n398, n409, n445);
  xor U311 ( n445, n406, n408);
  xor U312 ( n429, n461, n462);
  xor U313 ( n465, n467, n468);
  xor U314 ( n409, n417, n469);
  nand U315 ( n219, n224, n225);
  or U316 ( n221, n225, n224);
  xnor U317 ( n356, n357, n358);
  xnor U318 ( n399, n400, n401);
  xnor U319 ( n462, n463, n464);
  xnor U320 ( n265, n297, n275);
  xnor U321 ( n297, n276, n273);
  xnor U322 ( n289, n296, n333);
  xnor U323 ( n333, n293, n295);
  xnor U324 ( n441, n465, n466);
  xnor U325 ( n436, n455, n456);
  xnor U326 ( n455, n457, n458);
  xnor U327 ( n257, n250, n259);
  xnor U328 ( n259, n248, n251);
  xnor U329 ( n282, n265, n290);
  xnor U330 ( n290, n262, n264);
  nand U331 ( n295, n334, n335);
  or U332 ( n334, n319, n320);
  nand U333 ( n335, n321, n336);
  nand U334 ( n336, n320, n319);
  nand U335 ( n264, n291, n292);
  nand U336 ( n291, n296, n295);
  nand U337 ( n292, n293, n294);
  or U338 ( n294, n295, n296);
  nand U339 ( n251, n260, n261);
  nand U340 ( n260, n265, n264);
  nand U341 ( n261, n262, n263);
  or U342 ( n263, n264, n265);
  nand U343 ( n372, n419, n420);
  nand U344 ( n419, n398, n401);
  nand U345 ( n420, n400, n421);
  or U346 ( n421, n401, n398);
  nand U347 ( n281, n284, n285);
  nand U348 ( n284, n289, n288);
  nand U349 ( n285, n286, n287);
  or U350 ( n287, n288, n289);
  nand U351 ( n256, n277, n278);
  nand U352 ( n277, n282, n281);
  nand U353 ( n278, n279, n280);
  or U354 ( n280, n281, n282);
  nand U355 ( n236, n252, n253);
  nand U356 ( n252, n257, n256);
  nand U357 ( n253, n254, n255);
  or U358 ( n255, n256, n257);
  nand U359 ( n313, n374, n375);
  nand U360 ( n374, n355, n358);
  nand U361 ( n375, n357, n376);
  or U362 ( n376, n355, n358);
  and U363 ( n444, n449, n450);
  or U364 ( n449, n429, n430);
  nand U365 ( n450, n431, n451);
  nand U366 ( n451, n430, n429);
  nand U367 ( n358, n377, n378);
  or U368 ( n377, n341, n342);
  nand U369 ( n378, n343, n379);
  nand U370 ( n379, n342, n341);
  and U371 ( n230, n246, n247);
  nand U372 ( n246, n250, n251);
  nand U373 ( n247, n248, n249);
  or U374 ( n249, n250, n251);
  nand U375 ( n225, n232, n233);
  nand U376 ( n232, n237, n236);
  nand U377 ( n233, n234, n235);
  or U378 ( n235, n236, n237);
  and U379 ( n430, n452, n453);
  or U380 ( n452, n437, n438);
  nand U381 ( n453, n436, n454);
  nand U382 ( n454, n437, n438);
  nand U383 ( n401, n422, n423);
  nand U384 ( n422, n384, n385);
  nand U385 ( n423, n386, n424);
  or U386 ( n424, n385, n384);
  nand U387 ( n468, n473, n474);
  nand U388 ( n473, n461, n464);
  nand U389 ( n474, n463, n475);
  or U390 ( n475, n464, n461);
  nand U391 ( n464, n476, n477);
  nand U392 ( n476, n457, n456);
  nand U393 ( n477, n458, n478);
  or U394 ( n478, n456, n457);
  and U395 ( n276, n308, n309);
  nand U396 ( n308, n312, n313);
  nand U397 ( n309, n310, n311);
  or U398 ( n311, n312, n313);
  and U399 ( n408, n446, n447);
  or U400 ( n446, n441, n444);
  nand U401 ( n447, n443, n448);
  nand U402 ( n448, n444, n441);
  xnor U403 ( n361, n302, n299);
  xnor U404 ( n298, n267, n270);
  xnor U405 ( n469, n415, n418);
  xnor U406 ( n250, n244, n266);
  xnor U407 ( n266, n242, n245);
  xnor U408 ( n214, n351, n352);
  xnor U409 ( n351, n353, n354);
  xnor U410 ( n212, n329, n330);
  xnor U411 ( n329, n331, n332);
  xnor U412 ( n216, n394, n395);
  xnor U413 ( n394, n396, n397);
  xnor U414 ( n395, n435, n436);
  xnor U415 ( n435, n437, n438);
  xnor U416 ( n373, n367, n403);
  xnor U417 ( n403, n364, n366);
  xnor U418 ( n204, n318, n319);
  xnor U419 ( n318, n320, n321);
  xnor U420 ( n326, n340, n341);
  xnor U421 ( n340, n342, n343);
  xnor U422 ( n391, n428, n429);
  xnor U423 ( n428, n430, n431);
  xnor U424 ( n312, n360, n307);
  xnor U425 ( n360, n306, n267);
  nand U426 ( n288, n315, n316);
  nand U427 ( n315, n206, n205);
  nand U428 ( n316, n204, n317);
  or U429 ( n317, n205, n206);
  nand U430 ( n366, n404, n405);
  or U431 ( n404, n409, n408);
  nand U432 ( n405, n406, n407);
  nand U433 ( n407, n408, n409);
  and U434 ( n342, n380, n381);
  nand U435 ( n380, n350, n349);
  nand U436 ( n381, n348, n382);
  or U437 ( n382, n349, n350);
  and U438 ( n320, n337, n338);
  nand U439 ( n337, n328, n327);
  nand U440 ( n338, n326, n339);
  or U441 ( n339, n327, n328);
  and U442 ( n306, n368, n369);
  nand U443 ( n368, n373, n372);
  nand U444 ( n369, n370, n371);
  or U445 ( n371, n372, n373);
  and U446 ( n244, n271, n272);
  or U447 ( n271, n275, n276);
  nand U448 ( n272, n273, n274);
  nand U449 ( n274, n275, n276);
  nand U450 ( n349, n387, n388);
  or U451 ( n387, n353, n354);
  nand U452 ( n388, n352, n389);
  nand U453 ( n389, n353, n354);
  nand U454 ( n327, n344, n345);
  nand U455 ( n344, n331, n332);
  nand U456 ( n345, n330, n346);
  or U457 ( n346, n331, n332);
  nand U458 ( n205, n322, n323);
  or U459 ( n322, n209, n210);
  nand U460 ( n323, n208, n324);
  nand U461 ( n324, n209, n210);
  nand U462 ( n270, n299, n300);
  nand U463 ( n300, n301, n302);
  nand U464 ( n392, n432, n433);
  or U465 ( n432, n396, n397);
  nand U466 ( n433, n395, n434);
  nand U467 ( n434, n396, n397);
  and U468 ( n242, n267, n268);
  nand U469 ( n268, n269, n270);
  and U470 ( n417, n470, n471);
  nand U471 ( n470, n466, n468);
  nand U472 ( n471, n467, n472);
  or U473 ( n472, n468, n466);
  xnor U474 ( product_o[10], n289, n314);
  xnor U475 ( n314, n286, n288);
  nand U476 ( n229, n240, n241);
  or U477 ( n240, n245, n244);
  nand U478 ( n241, n242, n243);
  nand U479 ( n243, n244, n245);
  nand U480 ( n224, n226, n227);
  or U481 ( n226, n231, n230);
  nand U482 ( n227, n228, n229);
  nand U483 ( n228, n230, n231);
  nand U484 ( n385, n425, n426);
  nand U485 ( n425, n393, n392);
  nand U486 ( n426, n391, n427);
  or U487 ( n427, n392, n393);
  and U488 ( n301, n362, n363);
  nand U489 ( n362, n367, n366);
  nand U490 ( n363, n364, n365);
  or U491 ( n365, n366, n367);
  nand U492 ( n412, n413, n414);
  or U493 ( n413, n418, n417);
  nand U494 ( n414, n415, n416);
  nand U495 ( n416, n417, n418);
  and U496 ( n269, n303, n304);
  or U497 ( n303, n307, n306);
  nand U498 ( n304, n267, n305);
  nand U499 ( n305, n306, n307);
  xnor U500 ( product_o[8], n207, n208);
  xnor U501 ( n207, n209, n210);
  nand U502 ( n223, op2_i[7], op1_i[7]);
  nand U503 ( n222, n221, n219);
  and U504 ( n457, op2_i[2], n460, op1_i[2]);
  xnor U505 ( n460, n481, n482);
  nand U506 ( n481, op1_i[3], op2_i[1]);
  and U507 ( n482, op1_i[4], op2_i[0]);
  xnor U508 ( n456, n479, n480);
  nand U509 ( n479, op1_i[4], op2_i[1]);
  and U510 ( n480, op1_i[5], op2_i[0]);
  nand U511 ( product_o[15], n219, n220);
  nand U512 ( n220, op1_i[7], n221, op2_i[7]);
  xnor U513 ( n466, n485, n486);
  nand U514 ( n485, op1_i[6], op2_i[1]);
  and U515 ( n486, op1_i[7], op2_i[0]);
  xnor U516 ( n440, n459, n460);
  nand U517 ( n459, op1_i[2], op2_i[2]);
  xnor U518 ( n461, n483, n484);
  nand U519 ( n483, op1_i[5], op2_i[1]);
  and U520 ( n484, op1_i[6], op2_i[0]);
  xnor U521 ( n218, n439, n440);
  nand U522 ( n439, op1_i[1], op2_i[3]);
  nand U523 ( n209, op1_i[0], n212, op2_i[7]);
  nand U524 ( n353, op1_i[0], n216, op2_i[5]);
  nand U525 ( n437, op2_i[3], n440, op1_i[1]);
  nand U526 ( n396, op2_i[4], n218, op1_i[0]);
  nand U527 ( n418, op2_i[2], op1_i[6]);
  nand U528 ( n438, op2_i[3], op1_i[2]);
  nand U529 ( n397, op2_i[4], op1_i[1]);
  nand U530 ( n354, op2_i[5], op1_i[1]);
  nand U531 ( n302, op1_i[7], n412);
  and U532 ( n367, n302, n410);
  nand U533 ( n410, n202, n411);
  nand U534 ( n411, op2_i[2], op1_i[7]);
  not U535 ( n202, n412);
  and U536 ( n458, op1_i[3], op2_i[2]);
  and U537 ( n431, op2_i[3], op1_i[3]);
  and U538 ( n393, op2_i[4], op1_i[2]);
  and U539 ( n350, op2_i[5], op1_i[2]);
  and U540 ( n463, op1_i[4], op2_i[2]);
  and U541 ( n415, op2_i[1], op1_i[7]);
  and U542 ( n400, op2_i[4], op1_i[4]);
  and U543 ( n364, op2_i[3], op1_i[6]);
  and U544 ( n331, op2_i[6], op1_i[0], n214);
  and U545 ( n386, op2_i[4], op1_i[3]);
  and U546 ( n467, op1_i[5], op2_i[2]);
  and U547 ( n443, op2_i[3], op1_i[4]);
  and U548 ( n406, op2_i[3], op1_i[5]);
  and U549 ( n267, op2_i[4], op1_i[6]);
  nand U550 ( n245, op2_i[5], op1_i[7]);
  nand U551 ( n210, op2_i[7], op1_i[1]);
  and U552 ( n332, op2_i[6], op1_i[1]);
  and U553 ( n343, op2_i[5], op1_i[3]);
  and U554 ( n299, op2_i[3], op1_i[7]);
  and U555 ( n321, op2_i[6], op1_i[3]);
  and U556 ( n273, op2_i[5], op1_i[6]);
  and U557 ( n328, op2_i[6], op1_i[2]);
  and U558 ( n206, op2_i[7], op1_i[2]);
  and U559 ( n357, op2_i[5], op1_i[4]);
  and U560 ( n293, op2_i[6], op1_i[4]);
  and U561 ( n286, op2_i[7], op1_i[3]);
  and U562 ( n262, op2_i[6], op1_i[5]);
  and U563 ( n248, op2_i[6], op1_i[6]);
  xnor U564 ( product_o[6], n213, n214);
  nand U565 ( n213, op2_i[6], op1_i[0]);
  xnor U566 ( product_o[7], n211, n212);
  nand U567 ( n211, op2_i[7], op1_i[0]);
  and U568 ( n370, op2_i[4], op1_i[5]);
  and U569 ( n310, op2_i[5], op1_i[5]);
  xnor U570 ( product_o[5], n215, n216);
  nand U571 ( n215, op2_i[5], op1_i[0]);
  nand U572 ( n231, op2_i[6], op1_i[7]);
  xnor U573 ( product_o[4], n487, n218);
  nand U574 ( n487, op2_i[4], op1_i[0]);
  and U575 ( n279, op2_i[7], op1_i[4]);
  and U576 ( n254, op2_i[7], op1_i[5]);
  and U577 ( n234, op2_i[7], op1_i[6]);
  and U578 ( product_o[0], op2_i[0], op1_i[0]);
  and U579 ( product_o[1], op2_i[1], op1_i[0]);
  and U580 ( product_o[2], op2_i[2], op1_i[0]);
  and U581 ( product_o[3], op2_i[3], op1_i[0]);
endmodule
