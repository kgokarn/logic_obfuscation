module almost_correct_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493;

  xor U382 ( result_o[9], n262, n263);
  xor U383 ( n263, add2_i[9], add1_i[9]);
  xor U384 ( result_o[8], n268, n269);
  xor U385 ( n269, add2_i[8], add1_i[8]);
  xor U386 ( result_o[7], n273, n274);
  xor U387 ( n274, add2_i[7], add1_i[7]);
  xor U388 ( result_o[6], n286, n287);
  xor U389 ( n287, add2_i[6], add1_i[6]);
  xor U390 ( result_o[5], n290, n291);
  xor U391 ( n291, add2_i[5], add1_i[5]);
  xor U392 ( result_o[4], n294, n295);
  xor U393 ( n295, add2_i[4], add1_i[4]);
  xor U394 ( result_o[3], n298, n299);
  xor U395 ( n299, add2_i[3], add1_i[3]);
  xor U396 ( result_o[30], n316, n317);
  xor U397 ( result_o[2], n302, n321);
  xor U398 ( n321, add2_i[2], add1_i[2]);
  xor U399 ( result_o[29], n326, n327);
  xor U400 ( n327, add2_i[29], add1_i[29]);
  xor U401 ( result_o[28], n338, n339);
  xor U402 ( n339, add2_i[28], add1_i[28]);
  xor U403 ( result_o[27], n351, n352);
  xor U404 ( n352, add2_i[27], add1_i[27]);
  xor U405 ( result_o[26], n355, n356);
  xor U406 ( n356, add2_i[26], add1_i[26]);
  xor U407 ( result_o[25], n365, n366);
  xor U408 ( n366, add2_i[25], add1_i[25]);
  xor U409 ( result_o[24], n375, n376);
  xor U410 ( n376, add2_i[24], add1_i[24]);
  xor U411 ( result_o[23], n379, n380);
  xor U412 ( n380, add2_i[23], add1_i[23]);
  xor U413 ( result_o[22], n389, n390);
  xor U414 ( n390, add2_i[22], add1_i[22]);
  xor U415 ( result_o[21], n399, n400);
  xor U416 ( n400, add2_i[21], add1_i[21]);
  xor U417 ( result_o[20], n403, n404);
  xor U418 ( n404, add2_i[20], add1_i[20]);
  xor U419 ( result_o[1], n325, n413);
  xor U420 ( n413, add2_i[1], add1_i[1]);
  xor U421 ( result_o[19], n414, n415);
  xor U422 ( n415, add2_i[19], add1_i[19]);
  xor U423 ( result_o[18], n424, n425);
  xor U424 ( n425, add2_i[18], add1_i[18]);
  xor U425 ( result_o[17], n428, n429);
  xor U426 ( n429, add2_i[17], add1_i[17]);
  xor U427 ( result_o[16], n436, n437);
  xor U428 ( n437, add2_i[16], add1_i[16]);
  xor U429 ( result_o[15], n446, n447);
  xor U430 ( n447, add2_i[15], add1_i[15]);
  xor U431 ( result_o[14], n450, n451);
  xor U432 ( n451, add2_i[14], add1_i[14]);
  xor U433 ( result_o[13], n459, n460);
  xor U434 ( n460, add2_i[13], add1_i[13]);
  xor U435 ( result_o[12], n471, n472);
  xor U436 ( result_o[11], n479, n480);
  xor U437 ( result_o[10], n484, n485);
  xor U438 ( n485, add2_i[10], add1_i[10]);
  not U439 ( n228, n402);
  not U440 ( n223, n378);
  not U441 ( n218, n354);
  nor U442 ( n402, n398, n409);
  and U443 ( n409, n410, n394);
  nand U444 ( n410, n392, n411);
  nand U445 ( n411, n412, n406);
  nor U446 ( n378, n374, n385);
  and U447 ( n385, n386, n370);
  nand U448 ( n386, n368, n387);
  nand U449 ( n387, n388, n382);
  nor U450 ( n354, n350, n361);
  and U451 ( n361, n362, n344);
  nand U452 ( n362, n341, n363);
  nand U453 ( n363, n364, n358);
  nand U454 ( n340, n329, n220);
  not U455 ( n220, n341);
  not U456 ( n244, n478);
  not U457 ( n240, n439);
  not U458 ( n235, n417);
  not U459 ( n230, n392);
  not U460 ( n225, n368);
  not U461 ( n243, n462);
  not U462 ( n238, n449);
  not U463 ( n233, n427);
  nor U464 ( n350, n253, n219);
  nand U465 ( n290, n292, n293);
  nand U466 ( n293, n294, n285);
  nand U467 ( n349, n350, n342);
  nor U468 ( n454, n463, n464, n465);
  nor U469 ( n439, n435, n466);
  and U470 ( n466, n467, n241);
  nand U471 ( n467, n468, n469);
  or U472 ( n469, n470, n463);
  nor U473 ( n417, n412, n442);
  and U474 ( n442, n443, n407);
  nand U475 ( n443, n408, n444);
  nand U476 ( n444, n445, n440);
  nor U477 ( n392, n388, n420);
  and U478 ( n420, n421, n383);
  nand U479 ( n421, n384, n422);
  nand U480 ( n422, n423, n418);
  nor U481 ( n368, n364, n395);
  and U482 ( n395, n396, n359);
  nand U483 ( n396, n360, n397);
  nand U484 ( n397, n398, n393);
  nor U485 ( n341, n334, n371);
  and U486 ( n371, n372, n330);
  nand U487 ( n372, n332, n373);
  nand U488 ( n373, n374, n369);
  nor U489 ( n462, n458, n491);
  nor U490 ( n491, n489, n264);
  nor U491 ( n334, n254, n221);
  nor U492 ( n445, n261, n239);
  nor U493 ( n423, n259, n234);
  nor U494 ( n412, n260, n236);
  nor U495 ( n398, n257, n229);
  nor U496 ( n388, n258, n231);
  nor U497 ( n374, n255, n224);
  nor U498 ( n364, n256, n226);
  nor U499 ( n264, n453, n492);
  nor U500 ( n492, n270, n490);
  nor U501 ( n449, n445, n455);
  and U502 ( n455, n456, n441);
  nand U503 ( n456, n439, n457);
  nand U504 ( n457, n458, n454);
  nor U505 ( n427, n423, n432);
  and U506 ( n432, n433, n419);
  nand U507 ( n433, n417, n434);
  nand U508 ( n434, n435, n431);
  nand U509 ( n478, n266, n246, n245);
  nand U510 ( n441, n261, n239);
  nand U511 ( n419, n259, n234);
  nand U512 ( n394, n257, n229);
  nand U513 ( n370, n255, n224);
  nand U514 ( n344, n253, n219);
  nand U515 ( n407, n260, n236);
  nand U516 ( n383, n258, n231);
  nand U517 ( n359, n256, n226);
  nand U518 ( n330, n254, n221);
  nor U519 ( n318, n314, n320);
  nor U520 ( n474, n475, n476);
  nor U521 ( n475, n477, n465, n478);
  nor U522 ( n276, n278, n279);
  nand U523 ( n281, n483, n487);
  nand U524 ( n487, n283, n284, n250);
  not U525 ( n250, n292);
  nand U526 ( n476, n470, n482);
  or U527 ( n482, n462, n465);
  and U528 ( n320, n315, n333);
  nand U529 ( n333, n329, n331, n334);
  and U530 ( n277, n283, n284, n285);
  and U531 ( n431, n440, n407, n441);
  and U532 ( n406, n418, n383, n419);
  and U533 ( n382, n393, n359, n394);
  and U534 ( n358, n369, n330, n370);
  not U535 ( n251, n278);
  and U536 ( n329, n342, n343, n344);
  not U537 ( n245, n489);
  not U538 ( n246, n490);
  not U539 ( n242, n468);
  not U540 ( n241, n464);
  and U541 ( n483, n477, n488);
  nand U542 ( n488, n249, n284);
  not U543 ( n249, n288);
  not U544 ( n247, n272);
  not U545 ( n237, n408);
  not U546 ( n232, n384);
  not U547 ( n227, n360);
  not U548 ( n222, n332);
  not U549 ( n248, n267);
  nand U550 ( n306, n308, n309);
  nand U551 ( n308, add1_i[30], n311);
  nand U552 ( n309, add2_i[30], n310);
  or U553 ( n310, n311, add1_i[30]);
  or U554 ( n325, add2_i[0], add1_i[0]);
  or U555 ( n342, add2_i[26], add1_i[26]);
  nand U556 ( n286, n288, n289);
  nand U557 ( n289, n290, n283);
  nand U558 ( n337, n345, n346);
  nand U559 ( n345, add2_i[27], add1_i[27]);
  nand U560 ( n346, n347, n343);
  nand U561 ( n347, n348, n349);
  nand U562 ( n348, add2_i[26], add1_i[26]);
  nand U563 ( n294, n296, n297);
  nand U564 ( n296, add2_i[3], add1_i[3]);
  nand U565 ( n297, n298, n251);
  nand U566 ( n298, n300, n301);
  nand U567 ( n300, add2_i[2], add1_i[2]);
  nand U568 ( n301, n302, n252);
  not U569 ( n252, n279);
  nand U570 ( n302, n322, n323);
  nand U571 ( n322, add1_i[1], n325);
  nand U572 ( n323, add2_i[1], n324);
  or U573 ( n324, n325, add1_i[1]);
  not U574 ( n219, add1_i[25]);
  not U575 ( n253, add2_i[25]);
  xnor U576 ( result_o[31], n307, n306);
  xnor U577 ( n307, add1_i[31], add2_i[31]);
  and U578 ( n315, n335, n336);
  nand U579 ( n335, add2_i[28], add1_i[28]);
  nand U580 ( n336, n337, n331);
  nand U581 ( n311, n312, n313);
  nand U582 ( n312, add2_i[29], add1_i[29]);
  or U583 ( n313, n314, n315);
  nand U584 ( result_o[32], n303, n304);
  nand U585 ( n303, add1_i[31], n306);
  nand U586 ( n304, add2_i[31], n305);
  or U587 ( n305, n306, add1_i[31]);
  nor U588 ( n465, add2_i[10], add1_i[10]);
  nor U589 ( n463, add2_i[11], add1_i[11]);
  nor U590 ( n464, add2_i[12], add1_i[12]);
  nor U591 ( n278, add2_i[3], add1_i[3]);
  nor U592 ( n489, add2_i[9], add1_i[9]);
  nor U593 ( n279, add2_i[2], add1_i[2]);
  nor U594 ( n490, add2_i[8], add1_i[8]);
  nor U595 ( n267, n281, n282);
  and U596 ( n282, add1_i[3], n277, add2_i[3]);
  nor U597 ( n314, add2_i[29], add1_i[29]);
  nand U598 ( n408, add2_i[14], add1_i[14]);
  nand U599 ( n384, add2_i[17], add1_i[17]);
  nand U600 ( n360, add2_i[20], add1_i[20]);
  nand U601 ( n332, add2_i[23], add1_i[23]);
  or U602 ( n331, add2_i[28], add1_i[28]);
  or U603 ( n440, add2_i[14], add1_i[14]);
  or U604 ( n418, add2_i[17], add1_i[17]);
  or U605 ( n393, add2_i[20], add1_i[20]);
  or U606 ( n369, add2_i[23], add1_i[23]);
  or U607 ( n284, add2_i[6], add1_i[6]);
  or U608 ( n283, add2_i[5], add1_i[5]);
  or U609 ( n266, add2_i[7], add1_i[7]);
  nand U610 ( n484, n462, n486);
  nand U611 ( n486, n244, n281);
  nand U612 ( n446, n408, n448);
  nand U613 ( n448, n238, n440);
  nand U614 ( n424, n384, n426);
  nand U615 ( n426, n233, n418);
  nand U616 ( n414, n392, n416);
  nand U617 ( n416, n406, n235);
  nand U618 ( n399, n360, n401);
  nand U619 ( n401, n228, n393);
  nand U620 ( n389, n368, n391);
  nand U621 ( n391, n382, n230);
  nand U622 ( n375, n332, n377);
  nand U623 ( n377, n223, n369);
  nand U624 ( n365, n341, n367);
  nand U625 ( n367, n358, n225);
  nand U626 ( n351, n348, n353);
  nand U627 ( n353, n218, n342);
  nand U628 ( n338, n217, n340);
  not U629 ( n217, n337);
  nand U630 ( n262, n264, n265);
  nand U631 ( n265, n266, n246, n248);
  nand U632 ( n459, n439, n461);
  nand U633 ( n461, n454, n243);
  nand U634 ( n273, n247, n275);
  nand U635 ( n275, add2_i[1], add1_i[1], n276, n277);
  nand U636 ( n428, n427, n430);
  nand U637 ( n430, n242, n431, n241, n419);
  nand U638 ( n403, n402, n405);
  nand U639 ( n405, n237, n406, n407, n394);
  nand U640 ( n379, n378, n381);
  nand U641 ( n381, n232, n382, n383, n370);
  nand U642 ( n355, n354, n357);
  nand U643 ( n357, n227, n358, n359, n344);
  nand U644 ( n326, n320, n328);
  nand U645 ( n328, n222, n329, n330, n331);
  nand U646 ( n450, n449, n452);
  nand U647 ( n452, n453, n454, n245, n441);
  xnor U648 ( n479, add1_i[11], add2_i[11]);
  nor U649 ( n480, n481, n476);
  nor U650 ( n481, n478, n483, n465);
  xnor U651 ( n471, add1_i[12], add2_i[12]);
  nor U652 ( n472, n473, n242);
  nor U653 ( n473, n463, n474);
  xnor U654 ( n316, add1_i[30], add2_i[30]);
  nor U655 ( n317, n318, n319);
  and U656 ( n319, add1_i[29], add2_i[29]);
  nand U657 ( n272, n267, n280);
  nand U658 ( n280, add2_i[2], add1_i[2], n277, n251);
  nand U659 ( n270, add2_i[7], add1_i[7]);
  nand U660 ( n292, add2_i[4], add1_i[4]);
  nand U661 ( n288, add2_i[5], add1_i[5]);
  nand U662 ( n468, add2_i[11], add1_i[11]);
  and U663 ( n458, add1_i[9], add2_i[9]);
  and U664 ( n435, add2_i[12], add1_i[12]);
  or U665 ( n285, add2_i[4], add1_i[4]);
  and U666 ( n453, add2_i[8], add1_i[8]);
  or U667 ( n343, add2_i[27], add1_i[27]);
  nand U668 ( n477, add2_i[6], add1_i[6]);
  not U669 ( n239, add1_i[13]);
  not U670 ( n234, add1_i[16]);
  not U671 ( n236, add1_i[15]);
  not U672 ( n229, add1_i[19]);
  not U673 ( n231, add1_i[18]);
  not U674 ( n224, add1_i[22]);
  not U675 ( n226, add1_i[21]);
  not U676 ( n221, add1_i[24]);
  nand U677 ( n470, add2_i[10], add1_i[10]);
  not U678 ( n261, add2_i[13]);
  not U679 ( n259, add2_i[16]);
  not U680 ( n260, add2_i[15]);
  not U681 ( n257, add2_i[19]);
  not U682 ( n258, add2_i[18]);
  not U683 ( n255, add2_i[22]);
  not U684 ( n256, add2_i[21]);
  not U685 ( n254, add2_i[24]);
  nand U686 ( n436, n417, n438);
  nand U687 ( n438, n431, n240);
  nand U688 ( n268, n270, n271);
  nand U689 ( n271, n272, n266);
  nand U690 ( result_o[0], n325, n493);
  nand U691 ( n493, add2_i[0], add1_i[0]);
endmodule
