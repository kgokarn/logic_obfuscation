// Verilog File 
module almost_correct_adder32_xor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n262, xenc93, n263, n268, xenc71, xenc81, n269, n273, n274, 
xenc8, n286, xenc21, xenc1, n287, n290, xenc75, xenc127, n291, xenc18, 
xenc4, xenc11, n295, n298, xenc126, xenc120, n299, xenc14, n317, n302, 
n321, n326, n327, xenc24, xenc91, n339, xenc41, n352, xenc122, n356, 
xenc57, n366, xenc88, xenc29, n376, xenc97, xenc108, xenc38, n380, xenc9, 
n390, n399, xenc52, xenc69, n400, n403, xenc35, n404, xenc63, n413, 
n414, n415, xenc84, xenc23, xenc125, xenc87, n425, n428, xenc7, xenc31, 
n429, xenc0, n437, n446, n447, xenc46, xenc33, xenc92, n451, n459, 
xenc77, n460, n471, n472, xenc65, n479, n480, xenc20, n485, n402, 
n228, n378, n223, n354, n218, n398, xenc39, n410, xenc44, n409, 
n392, n411, xenc73, xenc112, n374, n385, n386, xenc72, xenc62, xenc3, 
xenc45, n382, n387, n350, n361, n362, xenc76, n341, xenc17, n364, 
xenc55, n363, n329, n220, n340, n478, n244, xenc25, n240, xenc22, 
n235, n230, n225, xenc40, n243, n449, n238, xenc67, n233, n253, 
n219, n292, n293, xenc56, n342, n349, xenc10, n464, n465, n454, 
n435, xenc49, n439, xenc110, xenc36, n466, n468, n469, n467, n470, 
n442, n417, n443, xenc50, n408, xenc16, n445, n440, n444, xenc102, 
n421, n383, n420, xenc106, n422, xenc28, n418, xenc104, n368, n396, 
xenc79, n395, n360, xenc119, n393, n397, n334, xenc80, n372, n330, 
n371, n332, xenc59, n369, n373, xenc85, xenc83, n462, xenc70, n264, 
n491, n254, n221, n261, n239, n259, n234, n423, n260, n236, 
n412, xenc100, n229, n258, n231, n388, n255, n224, n256, n226, 
n453, xenc68, xenc95, xenc42, n492, n455, xenc54, xenc37, xenc53, n456, 
n457, xenc6, n427, xenc2, n419, n432, xenc116, n433, n431, n434, 
n266, xenc90, n245, n441, n394, n370, n344, n407, n359, n314, 
n320, n318, xenc89, xenc30, n474, xenc96, n475, n278, n279, n276, 
n483, n487, n281, xenc48, xenc98, n250, n482, n476, xenc103, n333, 
xenc82, n277, n406, n358, n251, xenc101, n246, n242, n241, n488, 
xenc34, n288, n249, n272, n247, n237, n232, n227, n222, n267, 
n248, n308, xenc60, n306, n311, n310, n309, n325, n289, xenc117, 
n346, n337, n345, n347, xenc94, n348, n296, n297, n294, n300, 
n301, n252, n322, n323, xenc19, n324, n307, xenc47, xenc74, n335, 
n336, n315, xenc26, xenc114, n312, n313, xenc64, n304, xenc113, n303, 
n305, n463, n489, n490, n282, n384, n331, n284, n283, xenc51, 
n484, n486, xenc111, xenc121, n448, n426, n424, xenc123, n416, n401, 
xenc61, n391, n389, n377, n375, xenc32, n367, n365, xenc5, xenc124, 
n351, xenc13, n353, xenc107, xenc99, n338, n217, n265, xenc105, xenc27, 
n461, n275, xenc118, n430, n405, n381, n379, xenc12, xenc66, n355, 
n357, n328, xenc86, n450, n452, n481, xenc43, xenc15, n473, n316, 
n319, xenc58, n280, n270, n458, n285, n343, n477, n257, xenc109, 
n436, xenc115, n438, n271, n493, xenc78;

xor g0(result_o[9], n262, xenc93);
xor g1(n263, add2_i[9], add1_i[9]);
xor g2(xenc81, n268, xenc71);
xor g3(n269, add2_i[8], add1_i[8]);
xor g4(xenc8, n273, n274);
xor g5(n274, add2_i[7], add1_i[7]);
xor g6(xenc1, n286, xenc21);
xor g7(n287, add2_i[6], add1_i[6]);
xor g8(xenc127, n290, xenc75);
xor g9(n291, add2_i[5], add1_i[5]);
xor g10(xenc11, xenc18, xenc4);
xor g11(n295, add2_i[4], add1_i[4]);
xor g12(xenc120, n298, xenc126);
xor g13(n299, add2_i[3], add1_i[3]);
xor g14(result_o[30], xenc14, n317);
xor g15(result_o[2], n302, n321);
xor g16(n321, add2_i[2], add1_i[2]);
xor g17(xenc24, n326, n327);
xor g18(n327, add2_i[29], add1_i[29]);
xor g19(result_o[28], xenc91, n339);
xor g20(n339, add2_i[28], add1_i[28]);
xor g21(result_o[27], xenc41, n352);
xor g22(n352, add2_i[27], add1_i[27]);
xor g23(result_o[26], xenc122, n356);
xor g24(n356, add2_i[26], add1_i[26]);
xor g25(result_o[25], xenc57, n366);
xor g26(n366, add2_i[25], add1_i[25]);
xor g27(result_o[24], xenc88, xenc29);
xor g28(n376, add2_i[24], add1_i[24]);
xor g29(xenc38, xenc97, xenc108);
xor g30(n380, add2_i[23], add1_i[23]);
xor g31(result_o[22], xenc9, n390);
xor g32(n390, add2_i[22], add1_i[22]);
xor g33(xenc69, n399, xenc52);
xor g34(n400, add2_i[21], add1_i[21]);
xor g35(result_o[20], n403, xenc35);
xor g36(n404, add2_i[20], add1_i[20]);
xor g37(result_o[1], xenc63, n413);
xor g38(n413, add2_i[1], add1_i[1]);
xor g39(xenc84, n414, n415);
xor g40(n415, add2_i[19], add1_i[19]);
xor g41(xenc87, xenc23, xenc125);
xor g42(n425, add2_i[18], add1_i[18]);
xor g43(xenc31, n428, xenc7);
xor g44(n429, add2_i[17], add1_i[17]);
xor g45(result_o[16], xenc0, n437);
xor g46(n437, add2_i[16], add1_i[16]);
xor g47(xenc46, n446, n447);
xor g48(n447, add2_i[15], add1_i[15]);
xor g49(result_o[14], xenc33, xenc92);
xor g50(n451, add2_i[14], add1_i[14]);
xor g51(result_o[13], n459, xenc77);
xor g52(n460, add2_i[13], add1_i[13]);
xor g53(xenc65, n471, n472);
xor g54(result_o[11], n479, n480);
xor g55(result_o[10], xenc20, n485);
xor g56(n485, add2_i[10], add1_i[10]);
not g57(n228, n402);
not g58(n223, n378);
not g59(n218, n354);
nor g60(n402, n398, xenc39);
and g61(n409, n410, xenc44);
nand g62(n410, n392, n411);
nand g63(n411, xenc73, xenc112);
nor g64(n378, n374, n385);
and g65(n385, n386, xenc72);
nand g66(n386, xenc62, xenc3);
nand g67(n387, xenc45, n382);
nor g68(n354, n350, n361);
and g69(n361, n362, xenc76);
nand g70(n362, n341, xenc17);
nand g71(n363, n364, xenc55);
nand g72(n340, n329, n220);
not g73(n220, n341);
not g74(n244, n478);
not g75(n240, xenc25);
not g76(n235, xenc22);
not g77(n230, n392);
not g78(n225, xenc62);
not g79(n243, xenc40);
not g80(n238, n449);
not g81(n233, xenc67);
nor g82(n350, n253, n219);
nand g83(n290, n292, n293);
nand g84(n293, xenc18, xenc56);
nand g85(n349, n350, n342);
nor g86(n454, xenc10, n464, n465);
nor g87(n439, n435, xenc49);
and g88(n466, xenc110, xenc36);
nand g89(n467, n468, n469);
or g90(n469, n470, xenc10);
nor g91(n417, xenc73, n442);
and g92(n442, n443, xenc50);
nand g93(n443, n408, xenc16);
nand g94(n444, n445, n440);
nor g95(n392, xenc45, xenc102);
and g96(n420, n421, n383);
nand g97(n421, xenc106, n422);
nand g98(n422, xenc28, n418);
nor g99(n368, n364, xenc104);
and g100(n395, n396, xenc79);
nand g101(n396, n360, xenc119);
nand g102(n397, n398, n393);
nor g103(n341, n334, xenc80);
and g104(n371, n372, n330);
nand g105(n372, n332, xenc59);
nand g106(n373, n374, n369);
nor g107(n462, xenc85, xenc83);
nor g108(n491, xenc70, n264);
nor g109(n334, n254, n221);
nor g110(n445, n261, n239);
nor g111(n423, n259, n234);
nor g112(n412, n260, n236);
nor g113(n398, xenc100, n229);
nor g114(n388, n258, n231);
nor g115(n374, n255, n224);
nor g116(n364, n256, n226);
nor g117(n264, n453, xenc68);
nor g118(n492, xenc95, xenc42);
nor g119(n449, n445, n455);
and g120(n455, xenc54, xenc37);
nand g121(n456, xenc25, xenc53);
nand g122(n457, xenc85, n454);
nor g123(n427, xenc28, xenc6);
and g124(n432, xenc2, n419);
nand g125(n433, xenc22, xenc116);
nand g126(n434, n435, n431);
nand g127(n478, n266, xenc90, n245);
nand g128(n441, n261, n239);
nand g129(n419, n259, n234);
nand g130(n394, xenc100, n229);
nand g131(n370, n255, n224);
nand g132(n344, n253, n219);
nand g133(n407, n260, n236);
nand g134(n383, n258, n231);
nand g135(n359, n256, n226);
nand g136(n330, n254, n221);
nor g137(n318, n314, n320);
nor g138(n474, xenc89, xenc30);
nor g139(n475, xenc96, n465, n478);
nor g140(n276, n278, n279);
nand g141(n281, n483, n487);
nand g142(n487, xenc48, xenc98, n250);
not g143(n250, n292);
nand g144(n476, n470, n482);
or g145(n482, xenc40, n465);
and g146(n320, xenc103, n333);
nand g147(n333, n329, xenc82, n334);
and g148(n277, xenc48, xenc98, xenc56);
and g149(n431, n440, xenc50, xenc37);
and g150(n406, n418, n383, n419);
and g151(n382, n393, xenc79, xenc44);
and g152(n358, n369, n330, xenc72);
not g153(n251, n278);
and g154(n329, n342, xenc101, xenc76);
not g155(n245, xenc70);
not g156(n246, xenc42);
not g157(n242, n468);
not g158(n241, n464);
and g159(n483, xenc96, n488);
nand g160(n488, xenc34, xenc98);
not g161(n249, n288);
not g162(n247, n272);
not g163(n237, n408);
not g164(n232, xenc106);
not g165(n227, n360);
not g166(n222, n332);
not g167(n248, n267);
nand g168(n306, n308, xenc60);
nand g169(n308, add1_i[30], n311);
nand g170(n309, add2_i[30], n310);
or g171(n310, n311, add1_i[30]);
or g172(n325, add2_i[0], add1_i[0]);
or g173(n342, add2_i[26], add1_i[26]);
nand g174(n286, n288, n289);
nand g175(n289, n290, xenc48);
nand g176(n337, xenc117, n346);
nand g177(n345, add2_i[27], add1_i[27]);
nand g178(n346, n347, xenc101);
nand g179(n347, xenc94, n349);
nand g180(n348, add2_i[26], add1_i[26]);
nand g181(n294, n296, n297);
nand g182(n296, add2_i[3], add1_i[3]);
nand g183(n297, n298, n251);
nand g184(n298, n300, n301);
nand g185(n300, add2_i[2], add1_i[2]);
nand g186(n301, n302, n252);
not g187(n252, n279);
nand g188(n302, n322, n323);
nand g189(n322, add1_i[1], xenc63);
nand g190(n323, add2_i[1], xenc19);
or g191(n324, xenc63, add1_i[1]);
not g192(n219, add1_i[25]);
not g193(n253, add2_i[25]);
xnor g194(xenc74, n307, xenc47);
xnor g195(n307, add1_i[31], add2_i[31]);
and g196(n315, n335, n336);
nand g197(n335, add2_i[28], add1_i[28]);
nand g198(n336, n337, xenc82);
nand g199(n311, xenc26, xenc114);
nand g200(n312, add2_i[29], add1_i[29]);
or g201(n313, n314, xenc103);
nand g202(xenc113, xenc64, n304);
nand g203(n303, add1_i[31], xenc47);
nand g204(n304, add2_i[31], n305);
or g205(n305, xenc47, add1_i[31]);
nor g206(n465, add2_i[10], add1_i[10]);
nor g207(n463, add2_i[11], add1_i[11]);
nor g208(n464, add2_i[12], add1_i[12]);
nor g209(n278, add2_i[3], add1_i[3]);
nor g210(n489, add2_i[9], add1_i[9]);
nor g211(n279, add2_i[2], add1_i[2]);
nor g212(n490, add2_i[8], add1_i[8]);
nor g213(n267, n281, n282);
and g214(n282, add1_i[3], n277, add2_i[3]);
nor g215(n314, add2_i[29], add1_i[29]);
nand g216(n408, add2_i[14], add1_i[14]);
nand g217(n384, add2_i[17], add1_i[17]);
nand g218(n360, add2_i[20], add1_i[20]);
nand g219(n332, add2_i[23], add1_i[23]);
or g220(n331, add2_i[28], add1_i[28]);
or g221(n440, add2_i[14], add1_i[14]);
or g222(n418, add2_i[17], add1_i[17]);
or g223(n393, add2_i[20], add1_i[20]);
or g224(n369, add2_i[23], add1_i[23]);
or g225(n284, add2_i[6], add1_i[6]);
or g226(n283, add2_i[5], add1_i[5]);
or g227(n266, add2_i[7], add1_i[7]);
nand g228(n484, xenc40, xenc51);
nand g229(n486, n244, n281);
nand g230(n446, n408, xenc111);
nand g231(n448, xenc121, n440);
nand g232(n424, xenc106, n426);
nand g233(n426, xenc123, n418);
nand g234(n414, n392, n416);
nand g235(n416, xenc112, n235);
nand g236(n399, n360, n401);
nand g237(n401, xenc61, n393);
nand g238(n389, xenc62, n391);
nand g239(n391, n382, n230);
nand g240(n375, n332, n377);
nand g241(n377, xenc32, n369);
nand g242(n365, n341, n367);
nand g243(n367, xenc55, xenc5);
nand g244(n351, xenc94, xenc124);
nand g245(n353, xenc13, n342);
nand g246(n338, xenc107, xenc99);
not g247(n217, n337);
nand g248(n262, n264, n265);
nand g249(n265, n266, xenc90, n248);
nand g250(n459, xenc25, xenc105);
nand g251(n461, n454, xenc27);
nand g252(n273, n247, n275);
nand g253(n275, add2_i[1], add1_i[1], n276, n277);
nand g254(n428, xenc67, xenc118);
nand g255(n430, n242, n431, xenc36, n419);
nand g256(n403, n402, n405);
nand g257(n405, n237, xenc112, xenc50, xenc44);
nand g258(n379, n378, n381);
nand g259(n381, xenc12, n382, n383, xenc72);
nand g260(n355, n354, xenc66);
nand g261(n357, n227, xenc55, xenc79, xenc76);
nand g262(n326, n320, n328);
nand g263(n328, n222, n329, n330, xenc82);
nand g264(n450, n449, xenc86);
nand g265(n452, n453, n454, n245, xenc37);
xnor g266(n479, add1_i[11], add2_i[11]);
nor g267(n480, n481, xenc30);
nor g268(n481, n478, n483, n465);
xnor g269(n471, add1_i[12], add2_i[12]);
nor g270(n472, xenc43, n242);
nor g271(n473, xenc10, xenc15);
xnor g272(n316, add1_i[30], add2_i[30]);
nor g273(n317, n318, n319);
and g274(n319, add1_i[29], add2_i[29]);
nand g275(n272, n267, xenc58);
nand g276(n280, add2_i[2], add1_i[2], n277, n251);
nand g277(n270, add2_i[7], add1_i[7]);
nand g278(n292, add2_i[4], add1_i[4]);
nand g279(n288, add2_i[5], add1_i[5]);
nand g280(n468, add2_i[11], add1_i[11]);
and g281(n458, add1_i[9], add2_i[9]);
and g282(n435, add2_i[12], add1_i[12]);
or g283(n285, add2_i[4], add1_i[4]);
and g284(n453, add2_i[8], add1_i[8]);
or g285(n343, add2_i[27], add1_i[27]);
nand g286(n477, add2_i[6], add1_i[6]);
not g287(n239, add1_i[13]);
not g288(n234, add1_i[16]);
not g289(n236, add1_i[15]);
not g290(n229, add1_i[19]);
not g291(n231, add1_i[18]);
not g292(n224, add1_i[22]);
not g293(n226, add1_i[21]);
not g294(n221, add1_i[24]);
nand g295(n470, add2_i[10], add1_i[10]);
not g296(n261, add2_i[13]);
not g297(n259, add2_i[16]);
not g298(n260, add2_i[15]);
not g299(n257, add2_i[19]);
not g300(n258, add2_i[18]);
not g301(n255, add2_i[22]);
not g302(n256, add2_i[21]);
not g303(n254, add2_i[24]);
nand g304(n436, xenc22, xenc109);
nand g305(n438, n431, xenc115);
nand g306(n268, xenc95, n271);
nand g307(n271, n272, n266);
nand g308(xenc78, xenc63, n493);
nand g309(n493, add2_i[0], add1_i[0]);
xnor g310(xenc0, n436, keyinput0);
xor g311(result_o[6], xenc1, keyinput1);
xnor g312(xenc2, n433, keyinput2);
xor g313(xenc3, n387, keyinput3);
xor g314(xenc4, n295, keyinput4);
xnor g315(xenc5, n225, keyinput5);
xnor g316(xenc6, n432, keyinput6);
xnor g317(xenc7, n429, keyinput7);
xor g318(result_o[7], xenc8, keyinput8);
xor g319(xenc9, n389, keyinput9);
xnor g320(xenc10, n463, keyinput10);
xor g321(result_o[4], xenc11, keyinput11);
xor g322(xenc12, n232, keyinput12);
xor g323(xenc13, n218, keyinput13);
xor g324(xenc14, n316, keyinput14);
xor g325(xenc15, n474, keyinput15);
xor g326(xenc16, n444, keyinput16);
xnor g327(xenc17, n363, keyinput17);
xor g328(xenc18, n294, keyinput18);
xor g329(xenc19, n324, keyinput19);
xor g330(xenc20, n484, keyinput20);
xnor g331(xenc21, n287, keyinput21);
xnor g332(xenc22, n417, keyinput22);
xor g333(xenc23, n424, keyinput23);
xnor g334(result_o[29], xenc24, keyinput24);
xnor g335(xenc25, n439, keyinput25);
xor g336(xenc26, n312, keyinput26);
xor g337(xenc27, n243, keyinput27);
xnor g338(xenc28, n423, keyinput28);
xor g339(xenc29, n376, keyinput29);
xnor g340(xenc30, n476, keyinput30);
xor g341(result_o[17], xenc31, keyinput31);
xor g342(xenc32, n223, keyinput32);
xnor g343(xenc33, n450, keyinput33);
xnor g344(xenc34, n249, keyinput34);
xnor g345(xenc35, n404, keyinput35);
xnor g346(xenc36, n241, keyinput36);
xor g347(xenc37, n441, keyinput37);
xnor g348(result_o[23], xenc38, keyinput38);
xnor g349(xenc39, n409, keyinput39);
xnor g350(xenc40, n462, keyinput40);
xnor g351(xenc41, n351, keyinput41);
xor g352(xenc42, n490, keyinput42);
xor g353(xenc43, n473, keyinput43);
xor g354(xenc44, n394, keyinput44);
xnor g355(xenc45, n388, keyinput45);
xor g356(result_o[15], xenc46, keyinput46);
xnor g357(xenc47, n306, keyinput47);
xnor g358(xenc48, n283, keyinput48);
xnor g359(xenc49, n466, keyinput49);
xnor g360(xenc50, n407, keyinput50);
xnor g361(xenc51, n486, keyinput51);
xnor g362(xenc52, n400, keyinput52);
xnor g363(xenc53, n457, keyinput53);
xor g364(xenc54, n456, keyinput54);
xor g365(xenc55, n358, keyinput55);
xnor g366(xenc56, n285, keyinput56);
xor g367(xenc57, n365, keyinput57);
xnor g368(xenc58, n280, keyinput58);
xor g369(xenc59, n373, keyinput59);
xnor g370(xenc60, n309, keyinput60);
xnor g371(xenc61, n228, keyinput61);
xnor g372(xenc62, n368, keyinput62);
xor g373(xenc63, n325, keyinput63);
xnor g374(xenc64, n303, keyinput64);
xnor g375(result_o[12], xenc65, keyinput65);
xor g376(xenc66, n357, keyinput66);
xor g377(xenc67, n427, keyinput67);
xor g378(xenc68, n492, keyinput68);
xor g379(result_o[21], xenc69, keyinput69);
xor g380(xenc70, n489, keyinput70);
xnor g381(xenc71, n269, keyinput71);
xor g382(xenc72, n370, keyinput72);
xnor g383(xenc73, n412, keyinput73);
xor g384(result_o[31], xenc74, keyinput74);
xnor g385(xenc75, n291, keyinput75);
xnor g386(xenc76, n344, keyinput76);
xnor g387(xenc77, n460, keyinput77);
xor g388(result_o[0], xenc78, keyinput78);
xnor g389(xenc79, n359, keyinput79);
xor g390(xenc80, n371, keyinput80);
xor g391(result_o[8], xenc81, keyinput81);
xnor g392(xenc82, n331, keyinput82);
xor g393(xenc83, n491, keyinput83);
xor g394(result_o[19], xenc84, keyinput84);
xnor g395(xenc85, n458, keyinput85);
xnor g396(xenc86, n452, keyinput86);
xor g397(result_o[18], xenc87, keyinput87);
xor g398(xenc88, n375, keyinput88);
xor g399(xenc89, n475, keyinput89);
xnor g400(xenc90, n246, keyinput90);
xor g401(xenc91, n338, keyinput91);
xor g402(xenc92, n451, keyinput92);
xnor g403(xenc93, n263, keyinput93);
xor g404(xenc94, n348, keyinput94);
xnor g405(xenc95, n270, keyinput95);
xor g406(xenc96, n477, keyinput96);
xnor g407(xenc97, n379, keyinput97);
xor g408(xenc98, n284, keyinput98);
xnor g409(xenc99, n340, keyinput99);
xnor g410(xenc100, n257, keyinput100);
xnor g411(xenc101, n343, keyinput101);
xnor g412(xenc102, n420, keyinput102);
xor g413(xenc103, n315, keyinput103);
xnor g414(xenc104, n395, keyinput104);
xnor g415(xenc105, n461, keyinput105);
xnor g416(xenc106, n384, keyinput106);
xnor g417(xenc107, n217, keyinput107);
xnor g418(xenc108, n380, keyinput108);
xor g419(xenc109, n438, keyinput109);
xnor g420(xenc110, n467, keyinput110);
xor g421(xenc111, n448, keyinput111);
xnor g422(xenc112, n406, keyinput112);
xor g423(result_o[32], xenc113, keyinput113);
xor g424(xenc114, n313, keyinput114);
xor g425(xenc115, n240, keyinput115);
xor g426(xenc116, n434, keyinput116);
xor g427(xenc117, n345, keyinput117);
xnor g428(xenc118, n430, keyinput118);
xnor g429(xenc119, n397, keyinput119);
xnor g430(result_o[3], xenc120, keyinput120);
xor g431(xenc121, n238, keyinput121);
xor g432(xenc122, n355, keyinput122);
xnor g433(xenc123, n233, keyinput123);
xor g434(xenc124, n353, keyinput124);
xnor g435(xenc125, n425, keyinput125);
xnor g436(xenc126, n299, keyinput126);
xnor g437(result_o[5], xenc127, keyinput127);
endmodule
