library verilog;
use verilog.vl_types.all;
entity xnor_based_ripple_carry_adder32_tb is
end xnor_based_ripple_carry_adder32_tb;
