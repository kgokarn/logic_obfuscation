module xnor_based_carry_lookahead_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n412, n413, n414, n415, n417, n419, n421, n423, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n439,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n476, n477, n478, n479, n481, n482, n483, n484, n486, n487, n488,
         n489, n491, n492, n493, n494, n495, n496, n498, n499, n500, n501,
         n503, n504, n505, n506, n508, n509, n510, n511, n513, n514, n515,
         n516, n518, n519, n520, n521, n523, n524, n525, n526, n528, n529,
         n530, n531, n533, n534, n535, n536, n538, n539, n540, n541, n543,
         n544, n546, n547, n549, n550, n552, n553, n555, n556, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629;

  xor U464 ( result_o[9], n412, n413);
  xor U465 ( n413, add2_i[9], add1_i[9]);
  xor U466 ( result_o[8], n414, n415);
  xor U467 ( n415, add2_i[8], add1_i[8]);
  xor U473 ( result_o[31], n429, n430);
  xor U474 ( n430, add2_i[31], add1_i[31]);
  xor U475 ( result_o[30], n434, n435);
  xor U476 ( n435, add2_i[30], add1_i[30]);
  xor U478 ( result_o[29], n439, n442);
  xor U479 ( n442, add2_i[29], add1_i[29]);
  xor U480 ( result_o[28], n446, n447);
  xor U481 ( n447, add2_i[28], add1_i[28]);
  xor U482 ( result_o[27], n451, n452);
  xor U483 ( n452, add2_i[27], add1_i[27]);
  xor U484 ( result_o[26], n456, n457);
  xor U485 ( n457, add2_i[26], add1_i[26]);
  xor U486 ( result_o[25], n461, n462);
  xor U487 ( n462, add2_i[25], add1_i[25]);
  xor U488 ( result_o[24], n466, n467);
  xor U489 ( n467, add2_i[24], add1_i[24]);
  xor U490 ( result_o[23], n471, n472);
  xor U491 ( n472, add2_i[23], add1_i[23]);
  xor U492 ( result_o[22], n476, n477);
  xor U493 ( n477, add2_i[22], add1_i[22]);
  xor U494 ( result_o[21], n481, n482);
  xor U495 ( n482, add2_i[21], add1_i[21]);
  xor U496 ( result_o[20], n486, n487);
  xor U497 ( n487, add2_i[20], add1_i[20]);
  xor U498 ( n493, add2_i[1], add1_i[1]);
  xor U499 ( result_o[19], n491, n494);
  xor U500 ( n494, add2_i[19], add1_i[19]);
  xor U501 ( result_o[18], n498, n499);
  xor U502 ( n499, add2_i[18], add1_i[18]);
  xor U503 ( result_o[17], n503, n504);
  xor U504 ( n504, add2_i[17], add1_i[17]);
  xor U505 ( result_o[16], n508, n509);
  xor U506 ( n509, add2_i[16], add1_i[16]);
  xor U507 ( result_o[15], n513, n514);
  xor U508 ( n514, add2_i[15], add1_i[15]);
  xor U509 ( result_o[14], n518, n519);
  xor U510 ( n519, add2_i[14], add1_i[14]);
  xor U511 ( result_o[13], n523, n524);
  xor U512 ( n524, add2_i[13], add1_i[13]);
  xor U513 ( result_o[12], n528, n529);
  xor U514 ( n529, add2_i[12], add1_i[12]);
  xor U515 ( result_o[11], n533, n534);
  xor U516 ( n534, add2_i[11], add1_i[11]);
  xor U517 ( result_o[10], n538, n539);
  xor U518 ( n539, add2_i[10], add1_i[10]);
  not U519 ( n580, add2_i[7]);
  not U520 ( n586, add2_i[11]);
  not U521 ( n588, add2_i[20]);
  not U522 ( n582, add2_i[12]);
  nand U523 ( n496, add2_i[18], n568);
  or U524 ( n568, n498, add1_i[18]);
  not U525 ( n584, add2_i[21]);
  nand U526 ( n511, n569, add2_i[15]);
  or U527 ( n569, n513, add1_i[15]);
  or U528 ( n570, n581, n580);
  and U529 ( n617, n570, n571);
  and U530 ( n571, n572, n546);
  not U531 ( n572, add1_i[8]);
  or U532 ( n573, n587, n586);
  and U533 ( n583, n573, n574);
  and U534 ( n574, n575, n530);
  not U535 ( n575, add1_i[12]);
  or U536 ( n576, n589, n588);
  and U537 ( n585, n576, n577);
  and U538 ( n577, n578, n483);
  not U539 ( n578, add1_i[21]);
  or U540 ( n579, add2_i[0], add1_i[0]);
  not U541 ( n616, add2_i[8]);
  not U542 ( n608, add2_i[13]);
  or U543 ( n547, n580, n581);
  nor U544 ( n581, n417, add1_i[7]);
  or U545 ( n526, n582, n583);
  or U546 ( n479, n584, n585);
  not U547 ( n612, add2_i[5]);
  not U548 ( n626, add2_i[14]);
  not U549 ( n628, add2_i[29]);
  not U550 ( n614, add2_i[19]);
  not U551 ( n610, add2_i[22]);
  not U552 ( n618, add2_i[27]);
  not U553 ( n606, add2_i[10]);
  not U554 ( n624, add2_i[17]);
  or U555 ( n531, n586, n587);
  nor U556 ( n587, n533, add1_i[11]);
  or U557 ( n484, n588, n589);
  nor U558 ( n589, n486, add1_i[20]);
  not U559 ( n602, add2_i[6]);
  not U560 ( n604, add2_i[9]);
  not U561 ( n622, add2_i[16]);
  and U562 ( result_o[7], n417, n590);
  xnor U563 ( n590, add2_i[7], add1_i[7]);
  and U564 ( result_o[6], n419, n591);
  xnor U565 ( n591, add2_i[6], add1_i[6]);
  and U566 ( result_o[3], n425, n592);
  xnor U567 ( n592, add2_i[3], add1_i[3]);
  and U568 ( result_o[2], n441, n593);
  xnor U569 ( n593, add2_i[2], add1_i[2]);
  and U570 ( result_o[4], n423, n594);
  xnor U571 ( n594, add2_i[4], add1_i[4]);
  and U572 ( result_o[5], n421, n595);
  xnor U573 ( n595, add2_i[5], add1_i[5]);
  nor U574 ( n492, add2_i[0], add1_i[0]);
  not U575 ( n620, add2_i[4]);
  and U576 ( n607, n541, n596);
  and U577 ( n596, n540, n597);
  not U578 ( n597, add1_i[10]);
  or U579 ( n598, n623, n622);
  and U580 ( n625, n598, n599);
  and U581 ( n599, n600, n505);
  not U582 ( n600, add1_i[17]);
  or U583 ( n601, add2_i[0], add1_i[0]);
  nor U584 ( result_o[1], n492, n493);
  nand U585 ( n567, add2_i[0], add1_i[0]);
  or U586 ( n550, n603, n602);
  nor U587 ( n603, n419, add1_i[6]);
  or U588 ( n541, n605, n604);
  nor U589 ( n605, n412, add1_i[9]);
  or U590 ( n536, n606, n607);
  or U591 ( n521, n609, n608);
  nor U592 ( n609, n523, add1_i[13]);
  or U593 ( n474, n611, n610);
  nor U594 ( n611, n476, add1_i[22]);
  or U595 ( n553, n613, n612);
  nor U596 ( n613, n421, add1_i[5]);
  or U597 ( n489, n614, n615);
  nor U598 ( n615, n491, add1_i[19]);
  or U599 ( n544, n616, n617);
  or U600 ( n449, n618, n619);
  nor U601 ( n619, n451, add1_i[27]);
  or U602 ( n556, n620, n621);
  nor U603 ( n621, n423, add1_i[4]);
  or U604 ( n506, n622, n623);
  nor U605 ( n623, n508, add1_i[16]);
  or U606 ( n501, n624, n625);
  nand U607 ( n423, n558, n559);
  nand U608 ( n425, n561, n562);
  nand U609 ( n559, add2_i[3], n560);
  or U610 ( n516, n626, n627);
  nor U611 ( n627, n518, add1_i[14]);
  or U612 ( n437, n628, n629);
  nor U613 ( n629, n439, add1_i[29]);
  nand U614 ( n481, n483, n484);
  nand U615 ( n533, n536, n535);
  nand U616 ( n562, add2_i[2], n563);
  nand U617 ( n414, n546, n547);
  nand U618 ( n446, n449, n448);
  nand U619 ( result_o[0], n579, n567);
  nand U620 ( result_o[32], n426, n427);
  nand U621 ( n476, n478, n479);
  nand U622 ( n498, n501, n500);
  nand U623 ( n528, n530, n531);
  nand U624 ( n564, add1_i[1], n579);
  or U625 ( n566, n601, add1_i[1]);
  nand U626 ( n513, n515, n516);
  nand U627 ( n421, n556, n555);
  nand U628 ( n427, add2_i[31], n428);
  nand U629 ( n429, n431, n432);
  nand U630 ( n461, n463, n464);
  nand U631 ( n432, add2_i[30], n433);
  nand U632 ( n436, add1_i[29], n439);
  nand U633 ( n453, add1_i[26], n456);
  or U634 ( n455, n456, add1_i[26]);
  nand U635 ( n464, add2_i[24], n465);
  nand U636 ( n468, add1_i[23], n471);
  or U637 ( n470, n471, add1_i[23]);
  nand U638 ( n473, add1_i[22], n476);
  nand U639 ( n488, add1_i[19], n491);
  nand U640 ( n505, add1_i[16], n508);
  nand U641 ( n520, add1_i[13], n523);
  nand U642 ( n525, add1_i[12], n528);
  nand U643 ( n540, add1_i[9], n412);
  nand U644 ( n543, add1_i[8], n414);
  nand U645 ( n555, add1_i[4], n423);
  nand U646 ( n561, add1_i[2], n441);
  or U647 ( n563, n441, add1_i[2]);
  nand U648 ( n426, add1_i[31], n429);
  or U649 ( n428, n429, add1_i[31]);
  nand U650 ( n431, add1_i[30], n434);
  or U651 ( n433, n434, add1_i[30]);
  nand U652 ( n443, add1_i[28], n446);
  or U653 ( n445, n446, add1_i[28]);
  nand U654 ( n448, add1_i[27], n451);
  nand U655 ( n458, add1_i[25], n461);
  or U656 ( n460, n461, add1_i[25]);
  nand U657 ( n463, add1_i[24], n466);
  or U658 ( n465, n466, add1_i[24]);
  nand U659 ( n478, add1_i[21], n481);
  nand U660 ( n483, add1_i[20], n486);
  nand U661 ( n495, add1_i[18], n498);
  nand U662 ( n500, add1_i[17], n503);
  nand U663 ( n510, add1_i[15], n513);
  nand U664 ( n515, add1_i[14], n518);
  nand U665 ( n530, add1_i[11], n533);
  nand U666 ( n535, add1_i[10], n538);
  nand U667 ( n546, add1_i[7], n417);
  nand U668 ( n549, add1_i[6], n419);
  nand U669 ( n552, add1_i[5], n421);
  nand U670 ( n558, add1_i[3], n425);
  or U671 ( n560, n425, add1_i[3]);
  nand U672 ( n439, n443, n444);
  nand U673 ( n444, add2_i[28], n445);
  nand U674 ( n434, n436, n437);
  nand U675 ( n456, n458, n459);
  nand U676 ( n459, n460, add2_i[25]);
  nand U677 ( n451, n453, n454);
  nand U678 ( n454, add2_i[26], n455);
  nand U679 ( n471, n474, n473);
  nand U680 ( n466, n468, n469);
  nand U681 ( n469, n470, add2_i[23]);
  nand U682 ( n491, n495, n496);
  nand U683 ( n486, n489, n488);
  nand U684 ( n508, n510, n511);
  nand U685 ( n503, n505, n506);
  nand U686 ( n523, n525, n526);
  nand U687 ( n518, n521, n520);
  nand U688 ( n412, n544, n543);
  nand U689 ( n538, n541, n540);
  nand U690 ( n419, n553, n552);
  nand U691 ( n417, n550, n549);
  nand U692 ( n441, n565, n564);
  nand U693 ( n565, n566, add2_i[1]);
endmodule
