module ripple_carry_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107;

  xor U50 ( result_o[9], add2_i[9], n47);
  xor U51 ( result_o[8], add2_i[8], n48);
  xor U52 ( result_o[7], add2_i[7], n49);
  xor U53 ( result_o[6], add2_i[6], n50);
  xor U54 ( result_o[5], add2_i[5], n51);
  xor U55 ( result_o[4], add2_i[4], n52);
  xor U56 ( result_o[3], add2_i[3], n53);
  xor U57 ( result_o[2], add2_i[2], n54);
  xor U58 ( result_o[1], n55, add2_i[1]);
  xor U59 ( result_o[15], add2_i[15], n58);
  xor U60 ( n58, n59, add1_i[15]);
  xor U61 ( result_o[14], add2_i[14], n62);
  xor U62 ( n62, n63, add1_i[14]);
  xor U63 ( result_o[13], add2_i[13], n66);
  xor U64 ( n66, n67, add1_i[13]);
  xor U65 ( result_o[12], add2_i[12], n70);
  xor U66 ( n70, n71, add1_i[12]);
  xor U67 (  result_o[11], add2_i[11], n74);
  xor U68 ( n74, n75, add1_i[11]);
  xor U69 ( result_o[10], add2_i[10], n78);
  xor U70 ( n78, n79, add1_i[10]);
  xor U71 ( n47, n82, add1_i[9]);
  xor U72 ( n48, n85, add1_i[8]);
  xor U73 ( n49, n88, add1_i[7]);
  xor U74 ( n50, n91, add1_i[6]);
  xor U75 ( n51, n94, add1_i[5]);
  xor U76 ( n52, n97, add1_i[4]);
  xor U77 ( n53, n100, add1_i[3]);
  xor U78 ( n54, n103, add1_i[2]);
  xor U79 ( n55, n106, add1_i[1]);
  or U80 ( n106, add2_i[0], add1_i[0]);
  nand U81 ( n100, n101, n102);
  nand U82 ( n101, add1_i[2], n103);
  nand U83 ( n102, add2_i[2], n54);
  nand U84 ( n97, n98, n99);
  nand U85 ( n98, add1_i[3], n100);
  nand U86 ( n99, add2_i[3], n53);
  nand U87 ( n94, n95, n96);
  nand U88 ( n95, add1_i[4], n97);
  nand U89 ( n96, add2_i[4], n52);
  nand U90 ( n91, n92, n93);
  nand U91 ( n92, add1_i[5], n94);
  nand U92 ( n93, add2_i[5], n51);
  nand U93 ( n79, n80, n81);
  nand U94 ( n80, add1_i[9], n82);
  nand U95 ( n81, add2_i[9], n47);
  nand U96 ( n75, n76, n77);
  nand U97 ( n76, add1_i[10], n79);
  nand U98 ( n77, add2_i[10], n78);
  nand U99 ( n71, n72, n73);
  nand U100 ( n72, add1_i[11], n75);
  nand U101 ( n73, add2_i[11], n74);
  nand U102 ( n67, n68, n69);
  nand U103 ( n68, add1_i[12], n71);
  nand U104 ( n69, add2_i[12], n70);
  nand U105 ( n63, n64, n65);
  nand U106 ( n64, add1_i[13], n67);
  nand U107 ( n65, add2_i[13], n66);
  nand U108 ( n59, n60, n61);
  nand U109 ( n60, add1_i[14], n63);
  nand U110 ( n61, add2_i[14], n62);
  nand U111 ( n88, n89, n90);
  nand U112 ( n89, add1_i[6], n91);
  nand U113 ( n90, add2_i[6], n50);
  nand U114 ( n85, n86, n87);
  nand U115 ( n86, add1_i[7], n88);
  nand U116 ( n87, add2_i[7], n49);
  nand U117 ( n82, n83, n84);
  nand U118 ( n83, add1_i[8], n85);
  nand U119 ( n84, add2_i[8], n48);
  nand U120 ( n103, n104, n105);
  nand U121 ( n105, add1_i[1], n106);
  nand U122 ( n104, add2_i[1], n55);
  nand U123 ( result_o[16], n56, n57);
  nand U124 ( n56, add1_i[15], n59);
  nand U125 ( n57, add2_i[15], n58);
  nand U126 ( result_o[0], n106, n107);
  nand U127 ( n107, add2_i[0], add1_i[0]);
endmodule
