library verilog;
use verilog.vl_types.all;
entity array_multiplier8_tb is
end array_multiplier8_tb;
