library verilog;
use verilog.vl_types.all;
entity xnor_based_ripple_carry_adder16_tb is
end xnor_based_ripple_carry_adder16_tb;
