library verilog;
use verilog.vl_types.all;
entity underdesigned_multiplier8_tb is
end underdesigned_multiplier8_tb;
