library verilog;
use verilog.vl_types.all;
entity lower_part_or_ripple_carry_adder16_tb is
end lower_part_or_ripple_carry_adder16_tb;
