module ripple_carry_adder32 ( add1_i, add2_i, result_o );
  input [31:0] add1_i;
  input [31:0] add2_i;
  output [32:0] result_o;
  wire   n796, n797, n798, n799, n800, n801, n802, n803, n808, n809, n810,
         n811, n812, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n830, n831, n832, n833, n834,
         n835, n836, n837, n839, n840, n841, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n900, n901, n902, n903, n904, n905,
         n906, n907, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012;

  or U547 ( n886, add2_i[0], add1_i[0]);
  xor U562 ( result_o[8], n972, n812);
  xor U564 ( result_o[6], add2_i[6], n816);
  xor U565 ( result_o[5], add2_i[5], n817);
  xor U567 ( result_o[3], n819, n820);
  xor U568 ( n820, add2_i[3], add1_i[3]);
  xor U571 ( result_o[2], n837, add2_i[2]);
  xor U572 ( result_o[28], add2_i[28], n840);
  xor U573 ( result_o[27], add2_i[27], n846);
  xor U574 ( result_o[26], n856, n857);
  xor U575 ( result_o[25], n859, add2_i[25]);
  xor U577 ( result_o[24], n863, n864);
  xor U578 ( n864, add2_i[24], add1_i[24]);
  xor U579 ( result_o[23], add2_i[23], n867);
  xor U581 ( result_o[22], add2_i[22], n871);
  xor U583 ( result_o[21], add2_i[21], n875);
  xor U585 ( result_o[1], n886, n887);
  xor U586 ( n887, add2_i[1], add1_i[1]);
  xor U587 ( result_o[19], n884, add2_i[19]);
  xor U589 ( result_o[18], n894, n895);
  xor U590 ( result_o[15], add2_i[15], n907);
  xor U592 ( result_o[14], n912, n913);
  xor U593 ( n913, add2_i[14], add1_i[14]);
  xor U594 ( result_o[12], n921, add2_i[12]);
  xor U596 ( result_o[11], n926, n927);
  xor U597 ( n927, add2_i[11], add1_i[11]);
  xor U598 ( result_o[10], n930, add2_i[10]);
  xor U601 ( n837, n960, add1_i[2]);
  nand U602 ( n841, n796, n992);
  nand U603 ( n911, n1002, n915, n1001);
  nand U604 ( n995, n836, add2_i[28], add1_i[29], n998);
  xor U605 ( n977, n931, add1_i[10]);
  nand U606 ( n957, n965, n959, n958);
  not U607 ( n965, add1_i[3]);
  nand U608 ( n996, n841, add1_i[28], add1_i[29]);
  nand U609 ( n893, n800, n900, n901);
  nor U610 ( n974, n966, add1_i[11]);
  not U611 ( n966, n928);
  and U612 ( n985, n946, n988, n948);
  nor U613 ( n1000, n967, add1_i[24]);
  not U614 ( n967, n865);
  nand U615 ( n969, n902, add2_i[16], add1_i[17]);
  nand U616 ( n827, n976, n995, n996, n830);
  nand U617 ( n938, n937, n943, add2_i[6]);
  xor U618 ( n921, n922, add1_i[12]);
  xor U619 ( n871, n872, add1_i[22]);
  xor U620 ( n859, n855, add1_i[25]);
  nor U621 ( n840, n968, n981, n980);
  not U622 ( n968, n983);
  xnor U623 ( result_o[0], add2_i[0], add1_i[0]);
  xor U624 ( result_o[4], add2_i[4], n818);
  xnor U625 ( n903, n904, add1_i[16]);
  and U626 ( n896, add2_i[17], n893, n799);
  xnor U627 ( n880, n881, add1_i[20]);
  xor U628 ( result_o[31], n823, add2_i[31]);
  and U629 ( n848, n849, n850);
  not U630 ( n1003, add1_i[4]);
  nand U631 ( n897, n969, n970);
  or U632 ( n970, n800, n901);
  nand U633 ( n971, n909, n910);
  nand U634 ( n972, n815, n936);
  nand U635 ( n973, n977, add2_i[10]);
  nand U636 ( n925, n973, n974);
  nand U637 ( n975, n861, n860);
  not U638 ( n976, add1_i[30]);
  and U639 ( n815, n941, n942);
  and U640 ( n816, n943, n937);
  nand U641 ( n890, n892, n978);
  nor U642 ( n978, n897, add1_i[18]);
  and U643 ( n979, n817, n988);
  nor U644 ( n998, n980, n981);
  and U645 ( n980, add1_i[28], n990);
  and U646 ( n981, n991, add1_i[28]);
  or U647 ( n982, n991, add1_i[28], n990);
  or U648 ( n983, n991, add1_i[28], n990);
  or U649 ( n836, n991, add1_i[28], n990);
  nor U650 ( n984, n979, n986);
  nor U651 ( n937, n985, n986);
  nor U652 ( n986, n987, n946);
  not U653 ( n987, add1_i[6]);
  and U654 ( n988, add2_i[5], add1_i[6]);
  or U655 ( n989, n918, add1_i[13]);
  nor U656 ( n990, n992, n845);
  nor U657 ( n991, n797, n848);
  or U658 ( n916, n918, add1_i[13]);
  nor U659 ( n845, n797, n848);
  nand U660 ( n992, add2_i[27], n847);
  nand U661 ( n993, n909, n910);
  nand U662 ( n994, n933, n801, n934);
  and U663 ( n831, n995, n996);
  not U664 ( n997, add1_i[29]);
  nand U665 ( n999, n867, add2_i[23]);
  nand U666 ( n862, n999, n1000);
  nand U667 ( n1001, n989, add2_i[13]);
  not U668 ( n1002, add1_i[14]);
  xnor U669 ( n818, n954, n1003);
  not U670 ( n1005, add1_i[21]);
  not U671 ( n1004, add1_i[10]);
  xnor U672 ( n930, n931, n1004);
  xnor U673 ( n875, n876, n1005);
  not U674 ( n1006, add1_i[19]);
  not U675 ( n1007, add1_i[31]);
  xnor U676 ( n884, n885, n1006);
  xnor U677 ( n823, n824, n1007);
  not U678 ( n1012, add1_i[15]);
  not U679 ( n1011, add1_i[23]);
  nand U680 ( n830, n833, add2_i[29]);
  nand U681 ( n833, n834, n997, n835);
  nand U682 ( n850, add2_i[26], n851);
  nand U683 ( n851, n852, n798, n853);
  not U684 ( n801, add1_i[9]);
  xnor U685 ( n857, add2_i[26], n798);
  or U686 ( n948, n951, add1_i[5]);
  xor U687 ( result_o[30], n1008, n828);
  xor U688 ( n1008, add1_i[30], add2_i[30]);
  xor U689 ( result_o[29], n1009, n832);
  xor U690 ( n1009, add1_i[29], add2_i[29]);
  nand U691 ( n834, add1_i[28], n841);
  not U692 ( n802, add1_i[8]);
  xnor U693 ( result_o[20], add2_i[20], n880);
  nand U694 ( n933, add2_i[8], n939);
  nand U695 ( n940, add2_i[7], n944);
  nand U696 ( n852, add2_i[25], n854);
  nand U697 ( n945, add2_i[6], n943);
  not U698 ( n803, add1_i[7]);
  xnor U699 ( n894, add1_i[18], add2_i[18]);
  xnor U700 ( result_o[17], add2_i[17], n898);
  xnor U701 ( result_o[13], add2_i[13], n917);
  xnor U702 ( result_o[16], add2_i[16], n903);
  not U703 ( n800, add1_i[17]);
  xnor U704 ( n812, add2_i[8], n802);
  not U705 ( n798, add1_i[26]);
  xnor U706 ( result_o[7], add2_i[7], n1010);
  nand U707 ( n1010, n814, n815);
  xnor U708 ( result_o[9], add2_i[9], n808);
  not U709 ( n797, add1_i[27]);
  nand U710 ( n943, n946, n987, n947);
  nand U711 ( n885, n888, n889);
  xnor U712 ( n867, n868, n1011);
  xnor U713 ( n907, n993, n1012);
  or U714 ( n902, n904, add1_i[16]);
  or U715 ( n879, n881, add1_i[20]);
  nand U716 ( n917, n915, n989);
  nand U717 ( n910, n911, add2_i[14]);
  nand U718 ( n924, n925, add2_i[11]);
  nand U719 ( n922, n924, n923);
  nand U720 ( n855, n861, n860);
  nand U721 ( n861, add2_i[24], n862);
  nand U722 ( n947, n948, add2_i[5]);
  nand U723 ( n824, n825, n826);
  nand U724 ( n956, n957, add2_i[3]);
  nand U725 ( n914, n916, add2_i[13]);
  and U726 ( n846, n796, n847);
  nand U727 ( n826, n827, add2_i[30]);
  and U728 ( n817, n946, n948);
  nand U729 ( n958, add1_i[2], n960);
  nand U730 ( n954, n956, n955);
  nand U731 ( n952, add1_i[4], n954);
  nand U732 ( n847, n848, n797);
  nand U733 ( n873, add1_i[21], n876);
  nand U734 ( n889, n890, add2_i[18]);
  nand U735 ( n919, add1_i[12], n922);
  nand U736 ( n912, n914, n915);
  nand U737 ( n900, n902, add2_i[16]);
  nand U738 ( n960, n962, n961);
  nand U739 ( n962, n963, add2_i[1]);
  nand U740 ( n876, n877, n878);
  nand U741 ( n877, n879, add2_i[20]);
  nand U742 ( n821, add1_i[31], n824);
  nand U743 ( n863, n865, n866);
  nand U744 ( n865, n868, add1_i[23]);
  nand U745 ( n928, n931, add1_i[10]);
  nand U746 ( n931, n810, n932);
  nand U747 ( n939, n940, n802, n815);
  nand U748 ( n946, add1_i[5], n951);
  nand U749 ( n832, n834, n839);
  nand U750 ( n868, n870, n869);
  nand U751 ( n869, n872, add1_i[22]);
  nand U752 ( n905, n971, add1_i[15]);
  nand U753 ( n915, add1_i[13], n918);
  nand U754 ( n951, n953, n952);
  nand U755 ( n819, n959, n958);
  nand U756 ( n828, n831, n830);
  nand U757 ( n839, add2_i[28], n840);
  nand U758 ( n849, add1_i[26], n856);
  nand U759 ( n888, add1_i[18], n891);
  nand U760 ( n891, n892, n799);
  nand U761 ( n918, n919, n920);
  nand U762 ( n810, n935, add1_i[9]);
  nand U763 ( n934, add1_i[8], n811);
  nand U764 ( n898, n893, n799);
  nand U765 ( n835, add2_i[28], n982);
  nand U766 ( n856, n853, n858);
  nand U767 ( n853, add1_i[25], n975);
  or U768 ( n854, n975, add1_i[25]);
  nand U769 ( n872, n874, n873);
  nand U770 ( n878, add1_i[20], n881);
  nand U771 ( n892, add2_i[17], n893);
  nand U772 ( n926, n928, n929);
  nand U773 ( n935, n933, n934);
  nand U774 ( n809, n933, n801, n934);
  nand U775 ( n811, n815, n936);
  nand U776 ( result_o[32], n821, n822);
  nand U777 ( n808, n994, n810);
  nand U778 ( n860, add1_i[24], n863);
  nand U779 ( n881, n883, n882);
  nand U780 ( n883, add2_i[19], n884);
  nand U781 ( n901, add1_i[16], n904);
  nand U782 ( n904, n905, n906);
  nand U783 ( n923, add1_i[11], n926);
  nand U784 ( n932, add2_i[9], n809);
  nand U785 ( n936, add2_i[7], n814);
  nand U786 ( n955, add1_i[3], n819);
  nand U787 ( n961, add1_i[1], n886);
  or U788 ( n963, n886, add1_i[1]);
  nand U789 ( n822, add2_i[31], n823);
  nor U790 ( n895, n896, n897);
  nand U791 ( n825, add1_i[30], n828);
  not U792 ( n796, n991);
  nand U793 ( n858, n859, add2_i[25]);
  nand U794 ( n866, add2_i[23], n867);
  nand U795 ( n870, add2_i[22], n871);
  nand U796 ( n874, add2_i[21], n875);
  nand U797 ( n882, n885, add1_i[19]);
  not U798 ( n799, n897);
  nand U799 ( n906, add2_i[15], n907);
  nand U800 ( n909, add1_i[14], n912);
  nand U801 ( n920, add2_i[12], n921);
  nand U802 ( n929, add2_i[10], n930);
  nand U803 ( n944, n984, n803, n945);
  nand U804 ( n814, n984, n803, n938);
  nand U805 ( n942, add1_i[7], n816, add2_i[6]);
  or U806 ( n941, n984, n803);
  nand U807 ( n953, n818, add2_i[4]);
  nand U808 ( n959, add2_i[2], n837);
endmodule
