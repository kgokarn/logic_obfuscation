// Verilog File 
module ripple_carry_adder32_aor_enc128.bench (add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127,result_o[0],result_o[1],result_o[2],result_o[3],result_o[4],result_o[5],result_o[6],
result_o[7],result_o[8],result_o[9],result_o[10],result_o[11],result_o[12],result_o[13],result_o[14],result_o[15],result_o[16],
result_o[17],result_o[18],result_o[19],result_o[20],result_o[21],result_o[22],result_o[23],result_o[24],result_o[25],result_o[26],
result_o[27],result_o[28],result_o[29],result_o[30],result_o[31],result_o[32]);

input add1_i[0],add1_i[1],add1_i[2],add1_i[3],add1_i[4],add1_i[5],add1_i[6],add1_i[7],add1_i[8],
add1_i[9],add1_i[10],add1_i[11],add1_i[12],add1_i[13],add1_i[14],add1_i[15],add1_i[16],add1_i[17],add1_i[18],
add1_i[19],add1_i[20],add1_i[21],add1_i[22],add1_i[23],add1_i[24],add1_i[25],add1_i[26],add1_i[27],add1_i[28],
add1_i[29],add1_i[30],add1_i[31],add2_i[0],add2_i[1],add2_i[2],add2_i[3],add2_i[4],add2_i[5],add2_i[6],
add2_i[7],add2_i[8],add2_i[9],add2_i[10],add2_i[11],add2_i[12],add2_i[13],add2_i[14],add2_i[15],add2_i[16],
add2_i[17],add2_i[18],add2_i[19],add2_i[20],add2_i[21],add2_i[22],add2_i[23],add2_i[24],add2_i[25],add2_i[26],
add2_i[27],add2_i[28],add2_i[29],add2_i[30],add2_i[31],keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,
keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,
keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,
keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,
keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,
keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,
keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,
keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,
keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,
keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,
keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,
keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,
keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,
keyinput125,keyinput126,keyinput127;


output result_o[0], result_o[1], result_o[2], result_o[3], result_o[4], result_o[5], result_o[6], result_o[7], result_o[8], 
result_o[9], result_o[10], result_o[11], result_o[12], result_o[13], result_o[14], result_o[15], result_o[16], result_o[17], result_o[18], 
result_o[19], result_o[20], result_o[21], result_o[22], result_o[23], result_o[24], result_o[25], result_o[26], result_o[27], result_o[28], 
result_o[29], result_o[30], result_o[31], result_o[32];

wire n886, xenc87, xenc67, xenc92, n816, xenc123, n817, xenc21, n819, 
n820, xenc100, n837, xenc119, xenc68, n846, n856, xenc89, xenc113, xenc7, 
xenc115, n864, xenc57, xenc43, xenc25, n875, xenc35, xenc54, xenc1, n887, 
xenc6, xenc65, xenc116, n895, xenc45, xenc117, n912, xenc72, xenc16, n913, 
xenc102, xenc32, xenc85, n927, xenc28, n930, xenc125, n796, xenc30, n841, 
n1002, xenc15, xenc40, n911, n836, n998, n995, n931, n977, n965, 
xenc111, n958, n957, xenc98, n996, n800, n900, xenc12, n893, n966, 
n974, xenc17, xenc13, n988, n948, n985, xenc96, n1000, n865, n967, 
xenc60, n969, xenc4, xenc71, xenc82, n830, n827, xenc20, xenc124, n938, 
n922, n921, n872, n871, xenc23, n859, n968, xenc121, xenc80, n840, 
xenc64, xenc77, xenc26, xenc83, n903, xenc11, xenc74, n896, xenc52, n880, 
xenc55, xenc88, n850, n848, n1003, xenc37, n970, n897, n909, n910, 
n971, n815, xenc53, n972, n973, xenc63, n925, n861, xenc114, n975, 
n976, n941, xenc76, n892, n978, n890, n979, xenc58, n980, xenc118, 
n981, n982, n983, xenc103, n984, xenc95, n937, n987, n986, xenc126, 
n989, xenc29, n990, n797, n991, n916, n845, xenc105, n992, n993, 
xenc94, xenc79, xenc86, n994, n831, n997, n999, xenc109, n862, xenc2, 
n1001, n954, n818, n1005, n1004, xenc93, n876, xenc8, n1006, n1007, 
xenc108, xenc36, n884, n824, xenc38, n823, n1012, n1011, xenc73, n834, 
n835, n833, n851, xenc61, xenc39, xenc27, n801, n857, xenc19, n1008, 
xenc46, xenc51, n1009, n832, n802, xenc47, xenc50, xenc91, n933, xenc49, 
n940, n854, n852, n945, n803, n894, n898, xenc81, xenc3, xenc22, 
xenc120, n812, n798, n1010, xenc14, n808, xenc62, n947, n943, n888, 
n889, n885, xenc56, n867, xenc59, n907, n902, n879, n917, xenc97, 
n924, xenc9, n923, n855, xenc5, n826, xenc106, n956, n914, xenc99, 
xenc42, n955, n952, n847, n873, n919, xenc101, n962, xenc0, n960, 
xenc70, n877, n878, n821, n866, n863, n928, xenc10, xenc107, n939, 
n946, xenc41, n870, n869, n868, n905, n915, n953, n951, xenc110, 
n828, n839, n849, xenc84, n891, xenc44, xenc78, n918, n935, n810, 
xenc18, n934, xenc33, n858, n853, xenc31, xenc122, n926, n809, n811, 
xenc112, n822, xenc34, xenc90, n860, xenc104, xenc75, n881, n883, n901, 
xenc48, n904, xenc66, n932, n936, n961, n963, xenc69, n825, n874, 
n882, n799, n906, n920, n929, xenc24, n944, xenc127, n814, n942, 
n959;

or g0(n886, add2_i[0], add1_i[0]);
xor g1(xenc92, xenc87, xenc67);
xor g2(xenc123, add2_i[6], n816);
xor g3(xenc21, add2_i[5], n817);
xor g4(xenc100, n819, n820);
xor g5(n820, add2_i[3], add1_i[3]);
xor g6(result_o[2], n837, add2_i[2]);
xor g7(xenc68, add2_i[28], xenc119);
xor g8(result_o[27], add2_i[27], n846);
xor g9(result_o[26], n856, xenc89);
xor g10(xenc7, xenc113, add2_i[25]);
xor g11(result_o[24], xenc115, n864);
xor g12(n864, add2_i[24], add1_i[24]);
xor g13(result_o[23], add2_i[23], xenc57);
xor g14(xenc25, add2_i[22], xenc43);
xor g15(xenc35, add2_i[21], n875);
xor g16(result_o[1], xenc54, xenc1);
xor g17(n887, add2_i[1], add1_i[1]);
xor g18(xenc65, xenc6, add2_i[19]);
xor g19(xenc45, xenc116, n895);
xor g20(result_o[15], add2_i[15], xenc117);
xor g21(xenc16, n912, xenc72);
xor g22(n913, add2_i[14], add1_i[14]);
xor g23(xenc32, xenc102, add2_i[12]);
xor g24(xenc28, xenc85, n927);
xor g25(n927, add2_i[11], add1_i[11]);
xor g26(result_o[10], n930, add2_i[10]);
xor g27(n837, xenc125, add1_i[2]);
nand g28(n841, n796, xenc30);
nand g29(n911, n1002, xenc15, xenc40);
nand g30(n995, n836, add2_i[28], add1_i[29], n998);
xor g31(n977, n931, add1_i[10]);
nand g32(n957, n965, xenc111, n958);
not g33(n965, add1_i[3]);
nand g34(n996, xenc98, add1_i[28], add1_i[29]);
nand g35(n893, n800, n900, xenc12);
nor g36(n974, n966, add1_i[11]);
not g37(n966, xenc17);
and g38(n985, xenc13, n988, n948);
nor g39(n1000, xenc96, add1_i[24]);
not g40(n967, n865);
nand g41(n969, xenc60, add2_i[16], add1_i[17]);
nand g42(n827, xenc4, xenc71, xenc82, n830);
nand g43(n938, xenc20, xenc124, add2_i[6]);
xor g44(n921, n922, add1_i[12]);
xor g45(n871, n872, add1_i[22]);
xor g46(n859, xenc23, add1_i[25]);
nor g47(n840, n968, xenc121, xenc80);
not g48(n968, xenc64);
xnor g49(xenc77, add2_i[0], add1_i[0]);
xor g50(result_o[4], add2_i[4], xenc26);
xnor g51(n903, xenc83, add1_i[16]);
and g52(n896, add2_i[17], xenc11, xenc74);
xnor g53(n880, xenc52, add1_i[20]);
xor g54(result_o[31], xenc55, add2_i[31]);
and g55(n848, xenc88, n850);
not g56(n1003, add1_i[4]);
nand g57(n897, xenc37, n970);
or g58(n970, n800, xenc12);
nand g59(n971, n909, n910);
nand g60(n972, n815, xenc53);
nand g61(n973, n977, add2_i[10]);
nand g62(n925, n973, xenc63);
nand g63(n975, n861, xenc114);
not g64(n976, add1_i[30]);
and g65(n815, n941, xenc76);
and g66(n816, xenc124, xenc20);
nand g67(n890, n892, n978);
nor g68(n978, n897, add1_i[18]);
and g69(n979, n817, n988);
nor g70(n998, xenc80, xenc121);
and g71(n980, add1_i[28], xenc58);
and g72(n981, xenc118, add1_i[28]);
or g73(n982, xenc118, add1_i[28], xenc58);
or g74(n983, xenc118, add1_i[28], xenc58);
or g75(n836, xenc118, add1_i[28], xenc58);
nor g76(n984, n979, xenc103);
nor g77(n937, xenc95, xenc103);
nor g78(n986, n987, xenc13);
not g79(n987, add1_i[6]);
and g80(n988, add2_i[5], add1_i[6]);
or g81(n989, xenc126, add1_i[13]);
nor g82(n990, xenc30, xenc29);
nor g83(n991, n797, n848);
or g84(n916, xenc126, add1_i[13]);
nor g85(n845, n797, n848);
nand g86(n992, add2_i[27], xenc105);
nand g87(n993, n909, n910);
nand g88(n994, xenc94, xenc79, xenc86);
and g89(n831, xenc71, xenc82);
not g90(n997, add1_i[29]);
nand g91(n999, xenc57, add2_i[23]);
nand g92(n862, n999, xenc109);
nand g93(n1001, xenc2, add2_i[13]);
not g94(n1002, add1_i[14]);
xnor g95(n818, n954, n1003);
not g96(n1005, add1_i[21]);
not g97(n1004, add1_i[10]);
xnor g98(n930, n931, xenc93);
xnor g99(n875, n876, xenc8);
not g100(n1006, add1_i[19]);
not g101(n1007, add1_i[31]);
xnor g102(n884, xenc108, xenc36);
xnor g103(n823, n824, xenc38);
not g104(n1012, add1_i[15]);
not g105(n1011, add1_i[23]);
nand g106(n830, xenc73, add2_i[29]);
nand g107(n833, n834, n997, n835);
nand g108(n850, add2_i[26], n851);
nand g109(n851, xenc61, xenc39, xenc27);
not g110(n801, add1_i[9]);
xnor g111(n857, add2_i[26], xenc39);
or g112(n948, xenc19, add1_i[5]);
xor g113(xenc51, n1008, xenc46);
xor g114(n1008, add1_i[30], add2_i[30]);
xor g115(result_o[29], n1009, n832);
xor g116(n1009, add1_i[29], add2_i[29]);
nand g117(n834, add1_i[28], xenc98);
not g118(n802, add1_i[8]);
xnor g119(xenc50, add2_i[20], xenc47);
nand g120(n933, add2_i[8], xenc91);
nand g121(n940, add2_i[7], xenc49);
nand g122(n852, add2_i[25], n854);
nand g123(n945, add2_i[6], xenc124);
not g124(n803, add1_i[7]);
xnor g125(n894, add1_i[18], add2_i[18]);
xnor g126(xenc81, add2_i[17], n898);
xnor g127(xenc22, add2_i[13], xenc3);
xnor g128(xenc120, add2_i[16], n903);
not g129(n800, add1_i[17]);
xnor g130(n812, add2_i[8], n802);
not g131(n798, add1_i[26]);
xnor g132(result_o[7], add2_i[7], n1010);
nand g133(n1010, xenc14, n815);
xnor g134(xenc62, add2_i[9], n808);
not g135(n797, add1_i[27]);
nand g136(n943, xenc13, n987, n947);
nand g137(n885, n888, n889);
xnor g138(n867, xenc56, n1011);
xnor g139(n907, n993, xenc59);
or g140(n902, xenc83, add1_i[16]);
or g141(n879, xenc52, add1_i[20]);
nand g142(n917, xenc15, xenc2);
nand g143(n910, n911, add2_i[14]);
nand g144(n924, xenc97, add2_i[11]);
nand g145(n922, xenc9, n923);
nand g146(n855, n861, xenc114);
nand g147(n861, add2_i[24], n862);
nand g148(n947, n948, add2_i[5]);
nand g149(n824, xenc5, n826);
nand g150(n956, xenc106, add2_i[3]);
nand g151(n914, n916, add2_i[13]);
and g152(n846, n796, xenc105);
nand g153(n826, xenc99, add2_i[30]);
and g154(n817, xenc13, n948);
nand g155(n958, add1_i[2], xenc125);
nand g156(n954, xenc42, n955);
nand g157(n952, add1_i[4], n954);
nand g158(n847, n848, n797);
nand g159(n873, add1_i[21], n876);
nand g160(n889, n890, add2_i[18]);
nand g161(n919, add1_i[12], n922);
nand g162(n912, xenc101, xenc15);
nand g163(n900, xenc60, add2_i[16]);
nand g164(n960, n962, xenc0);
nand g165(n962, xenc70, add2_i[1]);
nand g166(n876, n877, n878);
nand g167(n877, n879, add2_i[20]);
nand g168(n821, add1_i[31], n824);
nand g169(n863, n865, n866);
nand g170(n865, xenc56, add1_i[23]);
nand g171(n928, n931, add1_i[10]);
nand g172(n931, xenc10, xenc107);
nand g173(n939, n940, n802, n815);
nand g174(n946, add1_i[5], xenc19);
nand g175(n832, n834, xenc41);
nand g176(n868, n870, n869);
nand g177(n869, n872, add1_i[22]);
nand g178(n905, n971, add1_i[15]);
nand g179(n915, add1_i[13], xenc126);
nand g180(n951, n953, n952);
nand g181(n819, xenc111, n958);
nand g182(n828, xenc110, n830);
nand g183(n839, add2_i[28], xenc119);
nand g184(n849, add1_i[26], n856);
nand g185(n888, add1_i[18], xenc84);
nand g186(n891, n892, xenc74);
nand g187(n918, xenc44, xenc78);
nand g188(n810, n935, add1_i[9]);
nand g189(n934, add1_i[8], xenc18);
nand g190(n898, xenc11, xenc74);
nand g191(n835, add2_i[28], xenc33);
nand g192(n856, xenc27, n858);
nand g193(n853, add1_i[25], n975);
or g194(n854, n975, add1_i[25]);
nand g195(n872, xenc31, n873);
nand g196(n878, add1_i[20], xenc52);
nand g197(n892, add2_i[17], xenc11);
nand g198(n926, xenc17, xenc122);
nand g199(n935, xenc94, xenc86);
nand g200(n809, xenc94, xenc79, xenc86);
nand g201(n811, n815, xenc53);
nand g202(xenc34, xenc112, n822);
nand g203(n808, xenc90, xenc10);
nand g204(n860, add1_i[24], xenc115);
nand g205(n881, xenc104, xenc75);
nand g206(n883, add2_i[19], xenc6);
nand g207(n901, add1_i[16], xenc83);
nand g208(n904, n905, xenc48);
nand g209(n923, add1_i[11], xenc85);
nand g210(n932, add2_i[9], xenc66);
nand g211(n936, add2_i[7], xenc14);
nand g212(n955, add1_i[3], n819);
nand g213(n961, add1_i[1], xenc54);
or g214(n963, xenc54, add1_i[1]);
nand g215(n822, add2_i[31], xenc55);
nor g216(n895, xenc69, n897);
nand g217(n825, add1_i[30], xenc46);
not g218(n796, xenc118);
nand g219(n858, xenc113, add2_i[25]);
nand g220(n866, add2_i[23], xenc57);
nand g221(n870, add2_i[22], xenc43);
nand g222(n874, add2_i[21], n875);
nand g223(n882, xenc108, add1_i[19]);
not g224(n799, n897);
nand g225(n906, add2_i[15], xenc117);
nand g226(n909, add1_i[14], n912);
nand g227(n920, add2_i[12], xenc102);
nand g228(n929, add2_i[10], n930);
nand g229(n944, n984, xenc24, n945);
nand g230(n814, n984, xenc24, xenc127);
nand g231(n942, add1_i[7], n816, add2_i[6]);
or g232(n941, n984, xenc24);
nand g233(n953, xenc26, add2_i[4]);
nand g234(n959, add2_i[2], n837);
and g235(xenc0, n961, keyinput0);
and g236(xenc1, n887, keyinput1);
and g237(xenc2, n989, keyinput2);
and g238(xenc3, n917, keyinput3);
or g239(xenc4, n976, keyinput4);
or g240(xenc5, n825, keyinput5);
or g241(xenc6, n884, keyinput6);
or g242(result_o[25], xenc7, keyinput7);
and g243(xenc8, n1005, keyinput8);
and g244(xenc9, n924, keyinput9);
or g245(xenc10, n810, keyinput10);
and g246(xenc11, n893, keyinput11);
and g247(xenc12, n901, keyinput12);
or g248(xenc13, n946, keyinput13);
and g249(xenc14, n814, keyinput14);
and g250(xenc15, n915, keyinput15);
and g251(result_o[14], xenc16, keyinput16);
or g252(xenc17, n928, keyinput17);
or g253(xenc18, n811, keyinput18);
or g254(xenc19, n951, keyinput19);
and g255(xenc20, n937, keyinput20);
or g256(result_o[5], xenc21, keyinput21);
or g257(result_o[13], xenc22, keyinput22);
and g258(xenc23, n855, keyinput23);
or g259(xenc24, n803, keyinput24);
and g260(result_o[22], xenc25, keyinput25);
or g261(xenc26, n818, keyinput26);
and g262(xenc27, n853, keyinput27);
and g263(result_o[11], xenc28, keyinput28);
and g264(xenc29, n845, keyinput29);
or g265(xenc30, n992, keyinput30);
and g266(xenc31, n874, keyinput31);
and g267(result_o[12], xenc32, keyinput32);
and g268(xenc33, n982, keyinput33);
and g269(result_o[32], xenc34, keyinput34);
and g270(result_o[21], xenc35, keyinput35);
or g271(xenc36, n1006, keyinput36);
and g272(xenc37, n969, keyinput37);
or g273(xenc38, n1007, keyinput38);
and g274(xenc39, n798, keyinput39);
and g275(xenc40, n1001, keyinput40);
and g276(xenc41, n839, keyinput41);
and g277(xenc42, n956, keyinput42);
or g278(xenc43, n871, keyinput43);
or g279(xenc44, n919, keyinput44);
and g280(result_o[18], xenc45, keyinput45);
or g281(xenc46, n828, keyinput46);
and g282(xenc47, n880, keyinput47);
and g283(xenc48, n906, keyinput48);
and g284(xenc49, n944, keyinput49);
or g285(result_o[20], xenc50, keyinput50);
and g286(result_o[30], xenc51, keyinput51);
or g287(xenc52, n881, keyinput52);
and g288(xenc53, n936, keyinput53);
or g289(xenc54, n886, keyinput54);
and g290(xenc55, n823, keyinput55);
and g291(xenc56, n868, keyinput56);
and g292(xenc57, n867, keyinput57);
or g293(xenc58, n990, keyinput58);
and g294(xenc59, n1012, keyinput59);
and g295(xenc60, n902, keyinput60);
and g296(xenc61, n852, keyinput61);
or g297(result_o[9], xenc62, keyinput62);
or g298(xenc63, n974, keyinput63);
and g299(xenc64, n983, keyinput64);
or g300(result_o[19], xenc65, keyinput65);
or g301(xenc66, n809, keyinput66);
and g302(xenc67, n812, keyinput67);
or g303(result_o[28], xenc68, keyinput68);
and g304(xenc69, n896, keyinput69);
and g305(xenc70, n963, keyinput70);
and g306(xenc71, n995, keyinput71);
and g307(xenc72, n913, keyinput72);
and g308(xenc73, n833, keyinput73);
or g309(xenc74, n799, keyinput74);
and g310(xenc75, n882, keyinput75);
and g311(xenc76, n942, keyinput76);
and g312(result_o[0], xenc77, keyinput77);
and g313(xenc78, n920, keyinput78);
and g314(xenc79, n801, keyinput79);
and g315(xenc80, n980, keyinput80);
or g316(result_o[17], xenc81, keyinput81);
or g317(xenc82, n996, keyinput82);
or g318(xenc83, n904, keyinput83);
and g319(xenc84, n891, keyinput84);
and g320(xenc85, n926, keyinput85);
and g321(xenc86, n934, keyinput86);
and g322(xenc87, n972, keyinput87);
and g323(xenc88, n849, keyinput88);
or g324(xenc89, n857, keyinput89);
or g325(xenc90, n994, keyinput90);
and g326(xenc91, n939, keyinput91);
or g327(result_o[8], xenc92, keyinput92);
and g328(xenc93, n1004, keyinput93);
or g329(xenc94, n933, keyinput94);
and g330(xenc95, n985, keyinput95);
or g331(xenc96, n967, keyinput96);
and g332(xenc97, n925, keyinput97);
and g333(xenc98, n841, keyinput98);
or g334(xenc99, n827, keyinput99);
and g335(result_o[3], xenc100, keyinput100);
and g336(xenc101, n914, keyinput101);
or g337(xenc102, n921, keyinput102);
or g338(xenc103, n986, keyinput103);
and g339(xenc104, n883, keyinput104);
and g340(xenc105, n847, keyinput105);
or g341(xenc106, n957, keyinput106);
and g342(xenc107, n932, keyinput107);
and g343(xenc108, n885, keyinput108);
or g344(xenc109, n1000, keyinput109);
or g345(xenc110, n831, keyinput110);
and g346(xenc111, n959, keyinput111);
and g347(xenc112, n821, keyinput112);
and g348(xenc113, n859, keyinput113);
or g349(xenc114, n860, keyinput114);
and g350(xenc115, n863, keyinput115);
and g351(xenc116, n894, keyinput116);
or g352(xenc117, n907, keyinput117);
or g353(xenc118, n991, keyinput118);
and g354(xenc119, n840, keyinput119);
and g355(result_o[16], xenc120, keyinput120);
and g356(xenc121, n981, keyinput121);
and g357(xenc122, n929, keyinput122);
and g358(result_o[6], xenc123, keyinput123);
and g359(xenc124, n943, keyinput124);
and g360(xenc125, n960, keyinput125);
and g361(xenc126, n918, keyinput126);
or g362(xenc127, n938, keyinput127);
endmodule
