module almost_correct_adder16 ( add1_i, add2_i, result_o );
  input [15:0] add1_i, add2_i;
  output [16:0] result_o;
  wire   n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202;

  xor U172 ( result_o[9], n98, n99);
  xor U173 ( n99, add2_i[9], add1_i[9]);
  xor U174 ( result_o[8], n106, n107);
  xor U175 ( n107, add2_i[8], add1_i[8]);
  xor U176 ( result_o[7], n115, n116);
  xor U177 ( n116, add2_i[7], add1_i[7]);
  xor U178 ( result_o[6], n119, n120);
  xor U179 ( n120, add2_i[6], add1_i[6]);
  xor U180 ( result_o[5], n131, n132);
  xor U181 ( n132, add2_i[5], add1_i[5]);
  xor U182 ( result_o[4], n134, n135);
  xor U183 ( n135, add2_i[4], add1_i[4]);
  xor U184 ( result_o[3], n138, n139);
  xor U185 ( n139, add2_i[3], add1_i[3]);
  xor U186 ( result_o[2], n142, n143);
  xor U187 ( n143, add2_i[2], add1_i[2]);
  xor U188 ( result_o[1], n147, n148);
  xor U189 ( n148, add2_i[1], add1_i[1]);
  xor U190 ( result_o[14], n162, n163);
  xor U191 ( n163, add2_i[14], add1_i[14]);
  xor U192 ( result_o[13], n166, n167);
  xor U193 ( n167, add2_i[13], add1_i[13]);
  xor U194 ( result_o[12], n178, n179);
  xor U195 ( n179, add2_i[12], add1_i[12]);
  xor U196 ( result_o[11], n189, n190);
  xor U197 ( n190, add2_i[11], add1_i[11]);
  xor U198 ( result_o[10], n195, n196);
  xor U199 ( n196, add2_i[10], add1_i[10]);
  not U200 ( n89, n100);
  not U201 ( n85, n165);
  nand U202 ( n157, n158, n159);
  nand U203 ( n159, n160, n161);
  nor U204 ( n102, n111, n200);
  nor U205 ( n127, n97, n95);
  nor U206 ( n183, n169, n201);
  nor U207 ( n201, n108, n200);
  nor U208 ( n100, n194, n198);
  and U209 ( n198, n102, n104, n127);
  nor U210 ( n165, n161, n173);
  and U211 ( n173, n170, n172, n88);
  not U212 ( n88, n174);
  and U213 ( n170, n184, n185);
  nand U214 ( n103, n97, n95);
  nand U215 ( n194, n183, n199);
  nand U216 ( n199, n92, n102);
  not U217 ( n92, n112);
  and U218 ( n122, n125, n103, n126);
  nand U219 ( n180, n170, n181);
  nand U220 ( n181, n174, n182);
  nand U221 ( n182, n171, n90);
  not U222 ( n90, n183);
  nand U223 ( n192, n174, n193);
  nand U224 ( n193, n171, n194);
  not U225 ( n93, n118);
  not U226 ( n96, n105);
  not U227 ( n91, n111);
  nand U228 ( n110, n112, n113);
  nand U229 ( n113, n94, n104);
  not U230 ( n94, n114);
  nand U231 ( n152, n154, n155);
  nand U232 ( n154, add1_i[14], n157);
  nand U233 ( n155, add2_i[14], n156);
  or U234 ( n156, n157, add1_i[14]);
  nand U235 ( n161, n175, n176);
  nand U236 ( n175, add2_i[12], add1_i[12]);
  nand U237 ( n176, n177, n172);
  nand U238 ( n188, add2_i[10], add1_i[10]);
  or U239 ( n185, add2_i[11], add1_i[11]);
  nand U240 ( n177, n186, n187);
  nand U241 ( n186, add2_i[11], add1_i[11]);
  nand U242 ( n187, n87, n185);
  not U243 ( n87, n188);
  nand U244 ( result_o[16], n149, n150);
  nand U245 ( n149, add1_i[15], n152);
  nand U246 ( n150, add2_i[15], n151);
  or U247 ( n151, n152, add1_i[15]);
  nor U248 ( n111, add2_i[7], add1_i[7]);
  nor U249 ( n200, add2_i[8], add1_i[8]);
  nor U250 ( n114, n127, n128);
  and U251 ( n128, n129, n103);
  nand U252 ( n129, n105, n130);
  nand U253 ( n130, add1_i[3], n125, add2_i[3]);
  or U254 ( n104, add2_i[6], add1_i[6]);
  nand U255 ( n174, add1_i[9], add2_i[9]);
  or U256 ( n171, add2_i[9], add1_i[9]);
  or U257 ( n147, add2_i[0], add1_i[0]);
  nand U258 ( n112, add2_i[6], add1_i[6]);
  nand U259 ( n105, add2_i[4], add1_i[4]);
  or U260 ( n172, add2_i[12], add1_i[12]);
  or U261 ( n125, add2_i[4], add1_i[4]);
  nand U262 ( n189, n188, n191);
  nand U263 ( n191, n192, n184);
  nand U264 ( n162, n158, n164);
  nand U265 ( n164, n85, n160);
  nand U266 ( n131, n105, n133);
  nand U267 ( n133, n134, n125);
  nand U268 ( n115, n112, n117);
  nand U269 ( n117, n118, n104);
  nand U270 ( n178, n86, n180);
  not U271 ( n86, n177);
  nand U272 ( n119, n93, n121);
  nand U273 ( n121, add2_i[1], add1_i[1], n122, n123);
  nand U274 ( n166, n165, n168);
  nand U275 ( n168, n169, n170, n171, n172);
  nand U276 ( n98, n100, n101);
  nand U277 ( n101, n96, n102, n103, n104);
  nand U278 ( n118, n114, n124);
  nand U279 ( n124, add1_i[2], n122, add2_i[2]);
  nand U280 ( n108, add2_i[7], add1_i[7]);
  nand U281 ( n158, add2_i[13], add1_i[13]);
  or U282 ( n123, add2_i[2], add1_i[2]);
  or U283 ( n126, add2_i[3], add1_i[3]);
  and U284 ( n169, add2_i[8], add1_i[8]);
  nand U285 ( n134, n136, n137);
  nand U286 ( n136, add2_i[3], add1_i[3]);
  nand U287 ( n137, n138, n126);
  nand U288 ( n138, n140, n141);
  nand U289 ( n140, add2_i[2], add1_i[2]);
  nand U290 ( n141, n142, n123);
  nand U291 ( n142, n144, n145);
  nand U292 ( n144, add1_i[1], n147);
  nand U293 ( n145, add2_i[1], n146);
  or U294 ( n146, n147, add1_i[1]);
  or U295 ( n160, add2_i[13], add1_i[13]);
  not U296 ( n95, add1_i[5]);
  not U297 ( n97, add2_i[5]);
  xnor U298 ( result_o[15], n153, n152);
  xnor U299 ( n153, add1_i[15], add2_i[15]);
  or U300 ( n184, add2_i[10], add1_i[10]);
  nand U301 ( n106, n108, n109);
  nand U302 ( n109, n110, n91);
  nand U303 ( n195, n174, n197);
  nand U304 ( n197, n171, n89);
  nand U305 ( result_o[0], n147, n202);
  nand U306 ( n202, add2_i[0], add1_i[0]);
endmodule
